�  �    9  X  x  �  �  �  �  �  	  D	  n	  �	  �	  �	  $
  V
  ~
  �
  �
    5  b  �  �  �  -  ^  �  �  �  '  X  �  �  �  -  b  �  �  �  1  h  �  �    7  r  �  �  
  <  ^  i  k  k  k  �  �    ,  K  j  �  �  �  �  �  	  D	  x	  �	  �	  �	  2
  s
  �
  �
  �
  .  e  �  �  �  .  Y  |  �  �  
  7  i  �  �    >  n  �  �    :  m  �  �  �  2  f  �  �  �  6  `  x  }  ~  �  �  �    &  C  a  �  �  �  �  	  N	  �	  �	  �	  

  8
  o
  �
  �
    6  Z  t  �  �  �    1  Y  �  �  �    O  }  �  �    J  {  �  �    C  v  �  �  	  <  r  �  �  
  .  =  A  A  A  '  �  �  "  I  d  �  �  �  #	  J	  y	  �	  �	  
  M
  {
  �
  �
  �
    $  Q  |  �  �  �  
  .  P  t  �  �  �     O  x  �  �    @  p  �  �     5  m  �  �    7  l  �  �  �    '  '  )  �  �  �    >  d  �  �  �  ;	  o	  �	  �	  �	  ;
  m
  �
  �
  �
  �
    .  L  l  �  �  �  �    $  P    �  �  �  )  Z  �  �  �    S  �  �  �    K  ~  �  �    F  y  �  �          �  +  �  �  0  \  �  �  	  <	  q	  �	  �	  	
  G
  {
  �
  �
  �
  �
  �
    7  Q  m  �  �  �  	  /  X  �  �  �  	  5  b  �  �  �    G  v  �  �  	  ;  n  �  �    5  g  �  �  �  	      S  �  �  �  .  ]  �  �  	  >	  p	  �	  �	  
  N
  `
  
  �
  �
  �
  �
    9  e  �  �  �  �    %  H  j  �  �  �    ?  h  �  �  �  &  Q  }  �  �    L  |  �  �    D  s  �  �        N  �  j  j  9  [  �  �  	  ?	  r	  �	  �	  
  J
  ^
  x
  �
  �
  �
  �
    3  O  o  �  �  �  �  �  $  R  �  �  �     /  `  �  �  �    K  ~  �  �    @  s  �  �    7  i  �  �        W  z  �  �  �  k  �  �  	  K	  ~	  �	  �	  %
  K
  j
  �
  �
  �
  �
  �
  �
    9  S  m  �  �  �    3  \  �  �  �    3  `  �  �  �    @  l  �  �  �  0  a  �  �  �  '  X  �  �  �       c  �  F  m  �  �  �  �  *	  ]	  �	  �	  �	  1
  >
  Z
  t
  �
  �
  �
  �
  �
    3  `  �  �  �  �      >  _    �  �  
  0  Y  �  �  �    C  m  �  �  	  8  k  �  �  �  2  a  �  �  �  *  �  �  O  o  �  	  	  
	  0	  ^	  �	  �	  �	  
  8
  Q
  f
  {
  �
  �
  �
    #  :  P  i  �  �  �  �  �    >  s  �  �  �     Q  �  �  �    4  o  �  �  �  /  a  �  �  �  %  V  �  �  �  $  �  �  l  `  o  �  �  "	  ;	  T	  l	  �	  �	  
  3
  ^
  q
  �
  �
  �
  �
  �
  �
    6  N  a  z  �  �     .  Q  x  �  �  
  5  b  �  �  �  #  P  �  �  �    L  y  �  �    ?  p  �  �  	  <  �  ^      T  r  �  �  4	  M	  n	  �	  �	  �	  6
  M
  [
  s
  �
  �
  �
  �
  �
  �
    G  |  �  �  �    N  �  �  �  �  -  \  �  �  �  "  T  �  �  �    D  v  �  �    >  q  �  �    7  h  �  �  �    !  L  }  �  �  :	  ^	  �	  �	  �	  
  3
  S
  h
  x
  �
  �
  �
    8  Y  x  �  �  	  5  ]  �  �  �    >  m  �  �    3  c  �  �  �  (  W  �  �  �     R  �  �  �    J  |  �    8  q  �    0  h  �  �  	  L	  j	  �	  �	  
  
  A
  }
  �
  �
  �
    >  n  �  �  �    E  r  �  �  �  *  Z  �  �  �    J  z  �  �    4  k  �  �  �  ,  ]  �  �  �  #  T  �  �  �  +  *  [  �    -  Z  o  �  �  1	  `	  �	  �	  �	  
  P
  �
  �
  �
    2  [  �  �  �    B  q  �  �  �  ,  [  �  �  �  '  U  �  �  �    L  |  �  �    E  v  �  �    =  n  �  �    ;  R  J    �  �  2  _  �  �  �  �  *	  U	  �	  �	  �	  
  O
  �
  �
  �
    K  {  �  �    9  k  �  �     .  [  �  �  �  '  S  �  �  �    P  �  �  �    I  |  �  �  
  =  q  �  �    6  �  �  �  �  �  �  �  .  t  �  �  �  0	  e	  �	  �	  �	  '
  W
  �
  �
  �
    O  �  �  �    D  v  �  �    =  m  �  �    4  c  �  �  �  0  `  �  �  �  )  ]  �  �  �  "  W  �  �  �    �  �  �  l  �  �  �    D  n  �  �  �  8	  r	  �	  �	  �	  %
  ]
  �
  �
  �
    N  �  �  �    >  q  �  �    5  g  �  �  �  /  `  �  �  �  (  X  �  �  �  %  V  �  �  �     S  �  �  �  �  �  i  �  �  �  �    7  T  �  �  �  	  =	  c	  �	  �	  �	  
  J
  x
  �
  �
    =  n  �  �  �  1  d  �  �  �  !  T  �  �  �    J  }  �  �    B  {  �  �    B  v  �  �    ?  q  �  ~  �  �  �  �  �  �    +  U  l  �  �  �  	  +	  R	  �	  �	  �	  
  4
  d
  �
  �
  �
  #  R  �  �  �    M  }  �  �    D  r  �  �    6  f  �  �  �  ,  _  �  �  �  /  e  �  �  �  -  a  t  �  �  �  �  �     C  X  a  �  �  �  �  �  �  !	  T	  �	  �	  �	  
  7
  i
  �
  �
  �
    N  �  �  �  
  <  o  �  �    8  i  �  �  �  /  _  �  �  �  &  V  �  �  �  !  V  �  �  �  $    �  �  �  �    (  P  f  t  �  �  �  �  �  	  -	  K	  j	  �	  �	  �	  
  B
  g
  �
  �
  �
    L  w  �  �  
  @  m  �  �  �  1  e  �  �  �  )  [  �  �  �    O  �  �  �    Q  �  �  �  �  �  �  �    '  9  X  v  �  �  �  �  �  	  +	  J	  f	  �	  �	  �	  �	  �	  
  5
  h
  �
  �
  �
  $  R  �  �  �    ?  r  �  �  	  9  j  �  �    3  c  �  �  �  .  ^  �  �  �  $  W  �  �  �  �  �    %  =  L  i  }  �  �  �  �  	  6	  K	  j	  �	  �	  �	  �	  �	  
  <
  \
  |
  �
  �
  �
    O  {  �  �  �  1  b  �  �  �     T  �  �  �    N  �  �  �    E  x  �  �    >  q  �  �  �  �    ,  G  T  j  �  �  �  �  �  	  4	  S	  w	  �	  �	  �	  
  
  <
  ]
  }
  �
  �
  �
    *  K  s  �  �    6  `  �  �  �  &  S  �  �  �    N  ~  �  �    J  {  �  �    D  u  �  �  �      <  X  l  �  �  �  �  �  
	  (	  G	  g	  �	  �	  �	  �	   
  !
  L
  �
  �
  �
  �
    4  Z  �  �  �  	  5  d  �  �  �    I  {  �  �  	  ;  n  �  �    4  f  �  �  �  0  a  �  �  �  �    #  D  `  u  �  �  �  �  	  !	  >	  [	  w	  �	  �	  �	  �	  

  1
  [
  �
  �
  �
  �
  /  b  �  �  �  	  8  g  �  �  �    K  z  �  �  	  :  m  �  �    4  f  �  �  �  0  ^  �  �  �  �  �    )  C  ]  q  �  �  �  �  	  0	  Q	  p	  �	  �	  �	  �	  
  ,
  P
  t
  �
  �
  �
    .  V  �  �  �    =  h  �  �  �  /  _  �  �  �  &  X  �  �  �  !  T  �  �  �    N  �  �  �  �  �      /  @  V  m  �  �  �  �  	  7	  [	  |	  �	  �	  �	  �	  
  C
  m
  �
  �
  �
  �
  "  E  n  �  �  �  #  Q  �  �  �    8  i  �  �  �  ,  _  �  �  �  (  Z  �  �  �  %  W  �  �  �  �  �    $  =  M  ^  |  �  �  �  �  	  <	  \	  }	  �	  �	  �	  �	  
  C
  r
  �
  �
  �
    A  n  �  �  �    @  n  �  �  �  "  R  �  �  �    L  �  �  �    J  |  �  �    E  r  �  �  �  �  �    #  B  Z  m  �  �  �  �  	  %	  E	  b	  �	  �	  �	  �	  �	  
  H
  r
  �
  �
  �
    D  n  �  �  �    F  q  �  �    6  e  �  �  �  /  b  �  �  �  .  a  �  �  �  ,  _  �  �  �  �  �  �       ?  W  h  y  �  �  �  �  (	  M	  l	  �	  �	  �	  �	  
  4
  Y
  �
  �
  �
  �
  !  E  f  �  �  �    D  u  �  �    9  l  �  �    >  q  �  �  
  =  p  �  �    ;  l  �  �  �  �  �  �       3  L  `  r  �  �  �  �  $	  N	  q	  �	  �	  �	  �	  
  3
  Y
  �
  �
  �
    /  Y    �  �  �  ,  ^  �  �  �  %  V  �  �  �  -  ]  �  �    8  h  �  �    ;  j  �  �  �  �  �  �  �  �    ,  E  ^  x  �  �  �  	  0	  P	  r	  �	  �	  �	  �	  
  2
  S
  �
  �
  �
    ,  b  �  �  �    K  �  �  �  #  R  �  �  �  +  \  �  �  �  1  c  �  �    8  n  �  �  �  �  �  �  �  �       =  V  n  �  �  �  �  	  6	  [	  y	  �	  �	  �	  
  ,
  N
  o
  �
  �
  �
    E  w  �  �    A  s  �  �    K  �  �  �  $  V  �  �  �  &  [  �  �  �  /  b  �  �  �            E  [  n    �  �  �  #  R  p  �  �  	  9	  g	  �	  �	  
  A
  s
  �
  �
     5  a  �  �  �  3  d  �  �  �  (  [  �  �  �  .  e  �  �  �  1  h  �  �    7  t  �  �    A  d  p  q  q  q  K  a  p  �  �  �    8  i  �  �  �  5	  k	  �	  �	  �	  .
  n
  �
  �
     7  m  �  �    <  v  �  �    6  m  �  �    E  y  �  �    A  t  �  �    H  �  �  �  !  S  �  �  �  �  �  �  X  g  |  �  �  �  +  `  �  �  �  -	  m	  �	  �	  �	  0
  k
  �
  �
    :  m  �  �    D  w  �  �    D  v  �  �  �  /  `  �  �  �  "  T  �  �  �    K  }  �  �    G  x  �  �  �  �  �  �  s  �  �  �  (  Z  �  �  �  	  Y	  �	  �	  �	   
  [
  �
  �
  �
  /  g  �  �    B  w  �  �  �    2  \  �  �  �    8  i  �  �  �  (  Y  �  �  �  ,  \  �  �  �  %  U  �  �  �  �  �    �  �  �  !  U  �  �  �  	  N	  �	  �	  �	  
  H
  �
  �
  �
  #  T  �  �  �  /  U  q  �  �  �  �  +  U    �  �    7  f  �  �  �  (  Z  �  �  �    Q  �  �  �    K  ~  �  �  �  �  A  �  �  �  $  L  x  �  �  *	  ]	  �	  �	  �	  0
  i
  �
  �
  �
  4  j  �  �       =  e  �  �  �    9  c  �  �  �    :  f  �  �  �  !  P  �  �  �    I  {  �  �    @  p  �  �  �  �  �  W  �  �    @  b  �  �  	  I	  x	  �	  �	  !
  Y
  �
  �
  �
  &  _  �  �  �  /  ]  |  �  �  �  �    @  n  �  �  �    J  {  �  �    0  e  �  �  �  -  ^  �  �  �  #  S  �  �  �  �  w  N  +  .    *  V  �  �  	  0	  Z	  �	  �	  
  9
  l
  �
  �
    @  }  �  �    B  _  w  �  �  �    7  _  �  �  �    B  r  �  �     2  d  �  �  �  (  [  �  �  �    R  �  �  �  �  �  �  O  o  3    6  b  �  �  	  ;	  f	  �	  �	  �	  >
  y
  �
  �
    O  �  �  �     ?  e  �  �  �    >  f  �  �  �    ;  g  �  �  �     M  ~  �  �    F  x  �  �    =  j  �  �  �  �  �  �  �  M  "  -  1  V  �  �  	  A	  o	  �	  �	  
  V
  �
  �
  �
  '  d  �  �     8  u  �  �  �  �    2  ]  �  �  �    <  m  �  �  �  !  P  �  �  �    N  �  �  �    D  u  �  �  �    w  �  .  g  m  M  R  �  �  	  ;	  f	  �	  �	  
  H
  {
  �
  �
    U  �  �  �  -  Y  v  �  �  �  �  $  R  v  �  �    1  ]  �  �  �    P  ~  �  �    C  v  �  �    :  p  �  �    �  �  �  �  �  I  \  U  s  �  �  	  P	  �	  �	  �	  )
  e
  �
  �
    C    �  �    +  L  |  �  �     '  W  �  �  �    :  j  �  �  �  -  `  �  �  �  '  X  �  �  �    P  �  �  �    �  W  e  �  �  (  ]  w  �  �  �  	  X	  �	  �	  �	  4
  m
  �
  �
  
  F    �  �    U  x  �  �  �  +  X  �  �  �    =  j  �  �  �  .  ^  �  �  �     P  �  �  �    M  �  �  �        .  z  u  �  �    \  ~  �  �  	  a	  �	  �	  �	  !
  \
  �
  �
  �
  +  e  �  �    7  n  �  �    E  w  �  �  
  =  l  �  �  �  -  _  �  �  �  !  Q  �  �  �    I  z  �  �    F  L  �  �  8  B  �  �    9  d  �  �  �  5	  o	  �	  �	  �	  0
  q
  �
  �
  �
  -  h  �  �    0  g  �  �    =  k  �  �    K  w  �  �    N  �  �  �    F  ~  �  �    ?  v  �  �    ;  I  r  �    4  e  �  �  �  9  b  �  �  �  5	  j	  �	  �	  �	  .
  g
  �
  �
  �
  *  ^  �  �  �  $  Y  �  �  �  !  S  �  �  �  %  P  �  �  �  $  S    �  �    S  �  �  �    L  �  �  �  t  �  �    *  f  �  �    >  f  �  �   	  ?	  j	  �	  �	  �	  -
  e
  �
  �
  �
     Y  �  �  �    O  �  �  �    I  }  �  �    I  {  �  �    I  x  �  �    G  w  �  �  
  ?  q  �  �  �  �  �    ,  a  h  �  �  !  Q  }  �  �  	  A	  n	  �	  �	  
  3
  a
  �
  �
  �
  %  X  �  �  �    O  �  �  �    G  z  �  �    A  u  �  �    ?  r  �  �  
  ;  n  �  �    6  f  �  �  �    �  	  (  V  �  �    '  Q  p  �  �  		  6	  b	  �	  �	  �	  )
  X
  �
  �
  �
    L  }  �  �    @  q  �  �  	  :  i  �  �    6  g  �  �  �  0  d  �  �  �  +  `  �  �  �  %  Z  �  �  �    H  W  z  �  �  �  �    =  q  �  �  �  !	  S	  �	  �	  �	  
  C
  v
  �
  �
  
  9  k  �  �  �  -  ]  �  �  �  !  R  �  �  �    K  }  �  �    N  ~  �  �    K  |  �  �    �  �    (  Q  p  T  m  z  �  �  �    >  e  �  �  �  '	  P	  v	  �	  �	  
  5
  b
  �
  �
  �
    Q  �  �  �    L    �  �    >  p  �  �    3  f  �  �     2  e  �  �    4  e  �  �  �    0  ;  P  S  w  z  �  �  �  �    )  Q  o  �  �  	  !	  B	  o	  �	  �	  �	  (
  T
  �
  �
  �
    D  t  �  �    @  q  �  �    :  i  �  �  �  -  ^  �  �  �  &  Z  �  �  �  %  Z  �    (  D  W  F  n    �  �  �  �    $  >  c  {  �  �  �  �  	  >	  q	  �	  �	  �	  #
  W
  �
  �
  �
    ?  t  �  �    6  h  �  �     /  `  �  �  �  %  U  �  �  �    T  �  �  �  "  V    %  <  P  U  m  �  �  �  �    #  >  Q  n  �  �  �  �  �  	  =	  ^	  �	  �	  �	  
  ;
  d
  �
  �
  �
    K  t  �  �    A  p  �  �    6  i  �  �  �  .  c  �  �  �  &  X  �  �  �  %  (  1  @  O  b  z  �  �  �  �    2  W  s  �  �  �  �  �  	  9	  X	  z	  �	  �	  �	  �	  
  <
  q
  �
  �
    -  \  �  �  �  !  Q  �  �  �    J    �  �    I  y  �  �    B  r  �  �    -  8  D  W  h  �  �  �  �       @  `  w  �  �  �  �  	  @	  ^	  {	  �	  �	  �	  �	  !
  L
  u
  �
  �
  �
    D  t  �  �  �  &  Z  �  �  �    L    �  �    E  x  �  �    @  r  �  �    2  :  K  [  v  �  �  �  �    .  G  d  z  �  �  �  �  	  I	  o	  �	  �	  �	  
  ,
  O
  t
  �
  �
  �
    <  d  �  �  �    F  p  �  �  
  9  i  �  �  �  1  a  �  �  �  *  ]  �  �  �    0  :  H  `  w  �  �  �    +  E  ]  z  �  �  �  �  	  5	  W	  |	  �	  �	  �	  
  *
  S
  �
  �
  �
    ;  e  �  �  �    I  w  �  �    6  e  �  �  �  .  `  �  �  �  *  \  �  �  �  �  �  .  9  F  a  �  �  �  �    5  T  o  �  �  �  �  	  0	  O	  n	  �	  �	  �	  �	  
  <
  e
  �
  �
  �
    @  r  �  �  �  &  X  �  �  �    N  �  �  �    I  |  �  �    G  x  �  �  �  �  �  /  ;  D  `  �  �  �  �    8  W  q  �  �  �  �  	  ;	  a	  	  �	  �	  �	  
  =
  b
  �
  �
  �
  �
  )  T  {  �  �    2  ^  �  �  �  )  Y  �  �  �  &  X  �  �  �  $  W  �  �  �        2  F  ]  |  �  �  �       >  X  s  �  �  �  �  	  @	  i	  �	  �	  �	  
  %
  E
  k
  �
  �
  �
    D  s  �  �    3  _  �  �  �  %  \  �  �  �  (  ]  �  �  �  %  [  �  �  �  �  �  �  �  8  H  W  k  �  �  �    7  S  m  �  �  �  �  
	  1	  U	  y	  �	  �	  �	  
  &
  G
  n
  �
  �
  �
    M  �  �  �    J  �  �  �    F  z  �  �    I  {  �  �    K  ~  �  �            3  >  M  e  �  �  �    <  ^    �  �  �  �  	  ?	  m	  �	  �	  �	  �	   
  E
  i
  �
  �
  �
    ?  t  �  �  
  9  l  �  �  
  B  t  �  �    D  v  �  �    F  x  �  �    .  7  7  7  7  2  <  N  g  �  �  �    <  ^  �  �  �  �  �  	  3	  j	  �	  �	  �	  

  A
  n
  �
  �
  �
  &  P    �  �    P  �  �  �    K  �  �  �    O  �  �  �  #  V  �  �  �  &  R  h  m  m  m  m  3  >  T  p  �  �    (  G  d  �  �  �  �  �   	  H	  {	  �	  �	  �	  1
  k
  �
  �
  �
     ]  �  �  �    R  �  �  �  $  X  �  �  �  *  [  �  �  �  /  h  �  �    :  l  �  �  �  �  �  �  =  I  e  �  �  �  �  +  K  d  �  �  �  	  ;	  d	  �	  �	  �	  #
  L
  y
  �
  �
    )  Z  �  �    -  \  �  �    5  k  �  �    B  s  �  �    D  w  �  �    S  �  �  �            �  �    9  \  �  �    >  f  �  �  	  8	  j	  �	  �	  
  @
  o
  �
  �
    D  s  �  �  
  F  w  �  �    ?  o  �  �    H  }  �  �    K  �  �  �    S  �  �  �  *  `  �  �  �  �  �  �  �    ;  j  �  �    R    �  �  #	  \	  �	  �	  �	  0
  i
  �
  �
  �
  :  p  �  �    @  y  �  �    @  v  �  �    N  �  �  �    N  �  �  �    V  �  �  �  .  a  �  �  �  %  ?  T  �  �    H  t  �  �  *  [  �  �  	  ?	  u	  �	  �	  	
  E
  {
  �
  �
    Q  �  �  �  )  ^  �  �    6  m  �  �    H  ~  �  �    Q  �  �  �  (  \  �  �  �  4  j  �  �    :  [  [  [  J  �     K  �  �     5  e  �  �  	  Q	  �	  �	  �	  )
  a
  �
  �
  �
  9  s  �  �    L  �  �  �  -  b  �  �    ;  q  �  �    U  �  �  �  2  f  �  �  �  1  e  �  �  �  '  R  ]  ]  _  p    (  P  �  �  
  ?  j  �  �  !	  T	  �	  �	  �	  3
  o
  �
  �
    F  �  �  �    [  �  �    9  q  �  �    Q  �  �  �  5  i  �  �    ;  l  �  �    2  b  �  �  �  ,  U  ]  `  `  �  �  <  ]  �  �    K  {  �  �  +	  `	  �	  �	  �	  7
  q
  �
  �
  	  E  �  �  �    W  �  �    6  n  �  �    K  �  �  �  ,  b  �  �    4  f  �  �  �  -  _  �  �  �  "  R  i  m  m    �  Y  s  �  �  )  S  �  �  �  8	  j	  �	  �	  
  R
  �
  �
  �
     \  �  �  �  0  k  �  �    B  ~  �  �  %  Z  �  �     0  _  �  �  �    N    �  �    E  w  �  �    :  k  w  w    �  �  �  �  �  $  Q  �  �  �  4	  j	  �	  �	  
  H
  
  �
  �
  $  ^  �  �  �  4  p  �  �    H  �  �  �  )  _  �  �  �  $  P  ~  �  �    G  w  �  �    >  n  �  �    8  k  v  v  '  V  �  �  �  �  #  C  n  �  �  	  N	  |	  �	  �	  )
  a
  �
  �
  �
  6  p  �  �    E  �  �  �  %  [  �  �  
  @  v  �  �    J  x  �  �  �  1  b  �  �  �  *  [  �  �  �    O  �  �  ?  v    Y  �       '  L  |  �  �  4	  d	  �	  �	  	
  H
  {
  �
  �
    V  �  �  �  .  j  �  �    F  �  �  �  ,  a  �  �  �    L  x  �  �    9  j  �  �  �  0  a  �  �  �  %  X  �  �  �    T  �  �    !  C  f  �  �  	  E	  x	  �	  �	  
  V
  �
  �
  �
  3  n  �  �    M  �  �  �  /  g  �  �    H  �  �  �    9  c  �  �  �  +  [  �  �  �  #  R  �  �  �    N  �  �  S  0  0  V  i  �    9  \  �  �  �  ,	  k	  �	  �	  

  F
  �
  �
  �
  '  a  �  �    B  {  �  �  '  ]  �  �  	  @  v  �  �    D  v  �  �    8  j  �  �  �  /  `  �  �  �  )  [  �  �  3  �  �  %  Y  �  �    8  k  �  �  &	  S	  	  �	  �	  -
  d
  �
  �
  �
  5  t  �  �    E  �  �  �    T  �  �  �  1  d  �  �    B  u  �  �    R  �  �  �  )  a  �  �  �  -  ]  �  i  �  �  �  �  /  [  �  �    >  o  �  �  %	  T	  	  �	  �	  )
  c
  �
  �
  �
  3  m  �  �    :  t  �  �    @  y  �  �    O  �  �  �  +  ]  �  �    7  j  �  �  	  ?  t  �  �    F  �    ]  �  �    M  �  �     (  M  �  �  �  6	  ]	  �	  �	  �	  1
  k
  �
  �
  �
  /  j  �  �  �  0  j  �  �    4  k  �  �  	  >  q  �  �    F  w  �  �    I  |  �  �    K  ~  �  �  �    I  �  �    3  G  �  �    ;  c  �  �  �  .	  ]	  �	  �	  �	  
  T
  �
  �
  �
    G  {  �  �    ?  t  �  �    4  l  �  �    4  b  �  �     1  a  �  �  �  -  ^  �  �  �  '  Z      f  �  �    4  c  �  �  �    7  o  �  �  �  .	  ^	  �	  �	  �	  (
  X
  �
  �
  �
  %  U  �  �  �    P  �  �  �    M  �  �  �    L  }  �  �    I  {  �  �    @  u  �  �  
  =  A  ^  �  �  �  �  �    J  z  �  �    =  g  �  �   	  5	  j	  �	  �	  �	  )
  ^
  �
  �
  �
     T  �  �  �    G  �  �  �    C  v  �  �    @  q  �  �    B  o  �  �    A  q  �  �    ~  �  �  +  l  v  �  �    ?  u  �  �    K  w  �  �   	  8	  h	  �	  �	  �	  +
  _
  �
  �
  �
    L  ~  �  �    B  v  �  �    ;  o  �  �    4  g  �  �    2  c  �  �  �  0  `  �  �  �  �  A  p  c  s  �  �  
  .  R  w  �  �    8  c  �  �  �  "	  N	  	  �	  �	  
  E
  t
  �
  �
    ;  i  �  �  �  ,  \  �  �  �  #  U  �  �  �    T  �  �  �    O  �  �  �    J    _  B  G  k  �  �  �  �  �    4  k  �  �  �  �  $  Z  �  �  �  	  9	  n	  �	  �	  �	  &
  X
  �
  �
  �
  "  R  �  �  �    G  w  �  �    :  k  �  �    4  j  �  �    ;  l  �  �    7  :  S  X  M  �  �  �      "  S  M  s  �  �  �  �  )  V  |  �  �  	  =	  j	  �	  �	  �	  "
  X
  �
  �
  �
    B  v  �  �  	  <  p  �  �     1  c  �  �  �  (  [  �  �  �  (  Y  �  �  �  ?  f  �  �  �  �  �    "  +  H  Z  x  �  �  �  �    1  Y    �  �  	  4	  Y	  �	  �	  �	  
  B
  o
  �
  �
    <  k  �  �    6  f  �  �  �  ,  ]  �  �  �    Q  �  �  �    T  �  �  4  G  �  �  �  �  �    2  F  [  y  �  �  �  �    %  F  g  }  �  �  �  �  )	  c	  �	  �	  �	  
  K
  �
  �
  �
    9  o  �  �    3  e  �  �  �  .  ]  �  �  �  *  Y  �  �  �  $  X  �  =  _  �  �  �  �     (  >  S  o  �  �  �  �    !  <  V  w  �  �  �  �  	  @	  f	  �	  �	  �	  
  D
  m
  �
  �
  �
  )  X  �  �  �    M  }  �  �    F  z  �  �  
  =  q  �  �    6  i  H  u  �  �  �  �  
    3  E  ]  w  �  �  �    >  ]  �  �  �  �  �  	  >	  `	  �	  �	  �	  �	  
  6
  b
  �
  �
  �
    I    �  �    E  t  �  �    >  q  �  �  
  <  m  �  �    7  h  x  �  �  �  �      *  J  d  �  �  �  �    $  G  d  �  �  �  �  	  <	  n	  �	  �	  �	  �	  
  E
  m
  �
  �
  �
    P  �  �  �  �  1  d  �  �  �  $  Z  �  �  �     R  �  �  �    O  z  �  �  �  �  �    3  C  [  }  �  �  �  �    4  R  m  �  �  �  �  	  ?	  k	  �	  �	  �	  
  P
  y
  �
  �
  �
  !  M  {  �  �    3  c  �  �  �  (  ]  �  �  �  '  Z  �  �  �  "  Q  V  V  �  �  �  �  �    0  A  P  f  �  �  �    .  K  p  �  �  �  �  	  8	  ]	  �	  �	  �	  �	  
  <
  `
  �
  �
  �
    J  |  �  �    H  w  �  �    M  }  �  �    K  |  �  �    E  [  [  [  �  �  �  �       +  A  S  p  �  �  �    ?  `  �  �  �  �  	  &	  V	  �	  �	  �	  �	  
  <
  b
  �
  �
  �
    C  z  �  �    7  o  �  �    9  m  �  �  	  :  l  �  �  	  ;  e  x  x  x  �  �  �      4  E  _  |  �  �  �    +  P  t  �  �  �  �  	  +	  _	  �	  �	  �	  
  =
  l
  �
  �
  �
    P  �  �  �    J  �  �  �  %  U  �  �  �  +  Y  �  �  �  1  ]  v  �  �  �  �  �  �  �    +  M  i    �  �  �     *  F  c  �  �  �  �  	  -	  T	  �	  �	  �	  �	  *
  a
  �
  �
  �
    S  �  �  �  '  [  �  �  �  .  `  �  �    6  f  �  �    <  q  �  �  �  �  �  �  �  �  �    -  L  e  x  �  �  �  �  "  I  h  �  �  �  ,	  M	  p	  �	  �	  �	  #
  J
  x
  �
  �
    B  u  �  �    =  u  �  �    H  |  �  �    M  ~  �  �    M    �  �            �  �  �    0  O  n  �  �  �  �    9  b  �  �  �  )	  W	  y	  �	  �	  
  B
  r
  �
  �
  	  @  o  �  �    =  l  �  �    8  i  �  �    9  t  �  �    ?  s  �  �    =  R  V  V  V  V  �  �  
  (  =  d  �  �  �  �  -  \  �  �  �  	  0	  e	  �	  �	  �	  !
  Z
  �
  �
  �
    X  �  �  �    M  �  �  �  $  W  �  �  �  %  W  �  �  �  &  a  �  �  �  .  b  �  �  �  �  �  �  �  �    .  K    �  �    3  e  �  �   	  (	  Y	  �	  �	  �	  "
  P
  �
  �
  �
    B  q  �  �    D  s  �  �    F    �  �  "  T  �  �  �     T  �  �  �  .  c  �  �  �    (  (  (  (  �  �    ,  ]  �  �  �    R  �  �  �  	  D	  |	  �	  �	  
  J
  �
  �
  �
  "  X  �  �  �  5  i  �  �    @  v  �  �    Q  �  �  �  '  Z  �  �  �  2  f  �  �    ?  t  �  �       +  �  �    (  X  �  �    @  m  �  �  	  F	  x	  �	  �	  
  C
  v
  �
  �
    H  {  �  �  "  V  �  �  �  )  \  �  �    <  o  �  �    C  w  �  �    P  �  �  �  *  _  �  �    4  d  �  �  �    &  F  �  �    @  e  �  �  	  X	  �	  �	  �	  #
  X
  �
  �
  �
  )  `  �  �  �  1  j  �  �    =  t  �  �    M  �  �  �  "  W  �  �  �  0  d  �  �  	  ?  s  �  �    H  }  �  �  �  �  &  K  �  �  �  3  d  �  �  	  A	  r	  �	  �	  
  S
  �
  �
  �
  $  a  �  �  �  5  q  �  �    J  �  �  �  )  a  �  �    F  }  �  �  %  [  �  �  �  7  n  �  �    G  ~  �  �  _  �  �    I  �  �  �    E  z  �  �  .	  ]	  �	  �	  �	  @
  u
  �
  �
    S  �  �  �  +  j  �  �    F  �  �  �  ,  a  �  �    H  ~  �  �  .  d  �  �    F  ~  �  �  $  `  �  �    �    �  �  "  Y  �  �     +  W  �  �  	  @	  o	  �	  �	  
  Q
  �
  �
  �
  &  d  �  �    8  u  �  �    O  �  �  �  3  h  �  �    L  ~  �  �  (  `  �  �    @  y  �  �    X  �  �  d  �  �  �     #  K  �  �    <  k  �  �  !	  T	  �	  �	  �	  .
  f
  �
  �
    >  z  �  �    T  �  �    7  n  �  �    O  �  �     8  n  �  �    T  �  �  �  3  m  �  �    N  �  �  W  5  4  J  �    L  �  �    1  Z  �  �  	  F	  t	  �	  �	  
  X
  �
  �
  �
  .  l  �  �    G  �  �  �  +  b  �  �    F  }  �  �  -  c  �  �    I  �  �  �  (  c  �  �    D    �  r  �  /  K  [    3  f  �  �    G  q  �  �  !	  Y	  �	  �	  �	  6
  q
  �
  �
    N  �  �  �  .  h  �  �    G  �  �  �  *  a  �  �    E  |  �  �  %  ]  �  �    ?  x  �  �  !  Z  �  �  �  �  �  >  #  0  O  v  �  �  +  c  �  �  	  H	  �	  �	  �	  +
  g
  �
  �
    H  �  �  �  )  c  �  �    F  �  �  �  *  b  �  �    I  �  �  �  /  h  �  �    K  �  �  �  -  g  �  �  �  U  �    >  S  t  �  �     <  n  �  �   	  [	  �	  �	  �	  :
  w
  �
  �
    T  �  �  �  0  m  �  �    K  �  �  �  .  e  �  �    L  �  �  �  0  h  �  �    L  �  �  �  ,  f  �  �  k  e  }  �  �  *  M  s  �  �  *  `  �  �  	  J	  ~	  �	  �	  0
  i
  �
  �
    I  �  �  �  #  ^  �  �    8  s  �  �    Q  �  �     5  k  �  �    P  �  �  �  1  i  �  �    K  �  �    #  M  z  �  �  $  `  �  �    7  k  �  �  	  G	  |	  �	  �	  
  Q
  �
  �
  �
  )  a  �  �    9  o  �  �    I  ~  �  �  $  Y  �  �  �  2  h  �  �  	  @  w  �  �    N  �  �  �  �  �      H  �  �  �  &  D  �  �  �  4  ]  �  �  	  A	  p	  �	  �	  
  N
  �
  �
  �
    S  �  �  �    U  �  �  �  -  a  �  �  	  <  o  �  �    J  }  �  �    T  �  �  �  %  \  �  @  �  �      b  �  �    2  V  �  �    B  g  �  �  	  I	  x	  �	  �	  
  M
  
  �
  �
  
  K  �  �  �    H  �  �  �    M  �  �  �  +  [  �  �  �  .  `  �  �  �  0  d  �  �  �  /    _  �  �    =  Z  �  �    0  l  �  �    ?  f  �  �  	  B	  o	  �	  �	  �	  =
  q
  �
  �
  �
  -  l  �  �  �  +  ^  �  �  �  &  Z  �  �  �  *  V  �  �  �  +  Y  �  �  �  (  Y  �  �     }  �  �  �  8  q  �  �    B  s  �  �    A  m  �  �  	  >	  m	  �	  �	  �	  6
  e
  �
  �
  �
  ,  a  �  �  �  #  X  �  �  �  !  T  �  �  �     P  �  �  �    O    �  �    K  |  �  Y  �  �  �  	  E  R  �  �  �  )  H  x  �  �    H  q  �  �  	  9	  i	  �	  �	  �	  0
  `
  �
  �
  �
  '  Z  �  �  �    Q  �  �  �    L  �  �  �    I  |  �  �    E  x  �  �    =  n  �  �  �  �  �    >  �  �  �    -  Q  �  �  �  
  7  j  �  �  �  /	  _	  �	  �	  �	  "
  S
  �
  �
  �
    F  y  �  �    =  o  �  �    ;  j  �  �    9  j  �  �    6  h  �  �  �  /  �  �  �  �  �  	  ?  u  �  �  �  �    G  p  �  �  �  /  a  �  �  �  	  N	  �	  �	  �	  
  A
  v
  �
  �
    2  d  �  �  �  &  Y  �  �  �    P  �  �  �     P  �  �  �    O    �  �  �  �  �  �    M    8  3  [  l  �  �    3  b  �  �  �  !  F  m  �  �  
	  4	  ]	  �	  �	  �	  %
  Z
  �
  �
  �
     R  �  �  �    D  t  �  �    8  j  �  �    5  m  �  �    5  j  �  �  �  �  �      "  ?  W    �  �  �  �    8  d  �  �  �    6  l  �  �  �  	  Q	  �	  �	  �	  
  >
  r
  �
  �
    =  n  �  �  	  7  e  �  �  �  ,  ^  �  �  �  (  Z  �  �  �  (  ^  �  �  �        1  A  ]  �  �  �  �  �  "  =  R  u  �  �  �  �  ;  n  �  �  �  	  U	  �	  �	  �	  
  =
  u
  �
  �
  �
  0  f  �  �  �  (  \  �  �  �    N  �  �  �    P  �  �  �  !  �  �  �  
    %  3  S  e  �  �  �  �    #  @  T  q  �  �  �  �  (  J  i  �  �  	  /	  Q	  x	  �	  �	  
  :
  e
  �
  �
    8  e  �  �  �  /  a  �  �  �  (  [  �  �  �    P  �  �  �  �  �  �        @  P  p  �  �  �    &  >  ]  {  �  �  �  �    8  a  ~  �  �  �   	  -	  e	  �	  �	  �	  
  L
  �
  �
  �
    =  r  �  �  	  <  m  �  �  
  7  f  �  �    3  c  �  �  �  �  �  
      N  ~  �  �  �  �    ;  X  z  �  �  �  �    9  X  w  �  �  �  	  -	  X	  {	  �	  �	  �	  2
  `
  �
  �
  �
    B  q  �  �     7  k  �  �  �  0  f  �  �  �  -  `  �  �      
    .  H  j  �  �  �  �       8  M  \  u  �  �  �  0  O  l  �  �  �  	  =	  `	  �	  �	  �	  �	  #
  F
  e
  �
  �
     &  S  �  �  �  $  Q  �  �  �  #  V  �  �  �  !  T  �  �  �          #  9  e  �  �  �    (  ?  X  u  �  �  �  �    >  f  �  �  �  �  	  2	  g	  �	  �	  �	  
  R
  �
  �
  �
    J  z  �  �    ?  o  �  �    B  s  �  �    @  s  �  �  �  �      
    -  L    �  �  �    ?  a    �  �  �  �  *  Q  o  �  �  �  �  	  2	  \	  �	  �	  �	  �	  3
  l
  �
  �
  �
  -  i  �  �  �  /  e  �  �    3  e  �  �  	  8  f  �  �  �  �  �        *  D  s  �  �  �    ,  N  p  �  �  �  �  �  1  Z  u  �  �  �  .	  U	  y	  �	  �	  �	  ,
  `
  �
  �
  �
  $  X  �  �  �    P  �  �  �    Q  �  �  �     R  �  �  �    "  "  "    +  <  O  d  �  �  �    '  B  k  �  �  �  �  �     T  ~  �  �  �  6	  a	  �	  �	  �	  '
  S
  �
  �
  �
    O  �  �  �    J  �  �  �    M  �  �  �    O  �  �  �  "  H  T  U  U  U  *  8  D  R  f  �  �  �    0  T  �  �  �    -  R    �  �  	  0	  _	  �	  �	  �	  
  <
  s
  �
  �
  �
  .  v  �  �    4  p  �  �  
  :  o  �  �    @  r  �  �    F  v  �  �  �  �  �  ;  B  K  c  �  �  �    7  T  v  �  �    <  f  �  �  	  ?	  c	  �	  �	  �	  
  A
  p
  �
  �
    ;  l  �  �    6  m  �  �    B  w  �  �    D  x  �  �    L  ~  �  �  �  �  �  �  �  G  ]  o  �  �  �    ;  g  �  �  �  +  W  �  �  �  !	  S	  �	  �	  �	  
  I
  }
  �
  �
    L  x  �  �    G  v  �  �    @  r  �  �    ?  z  �  �    C  y  �  �    G  `  c  c  c  c  Z  }  �  �  �  !  P  r  �  �    F  w  �  �  	  5	  g	  �	  �	  �	  .
  g
  �
  �
  �
  /  j  �  �  �  -  _  �  �  	  6  h  �  �    3  d  �  �    2  n  �  �  	  :  m  �  �  �  �  �  �  }  �  �    ;  ^  �  �  �    H  u  �  �  	  A	  x	  �	  �	  
  F
  {
  �
  �
    K    �  �  )  \  �  �  �  )  b  �  �    8  m  �  �    8  m  �  �  	  F  {  �  �    F  v          /  d  �  �    <  l  �  �  "  Q  �  �  
	  A	  s	  �	  �	  
  U
  �
  �
  �
  )  d  �  �    <  u  �  �    O  �  �  �  /  d  �  �    D  y  �  �    T  �  �  �  ,  b  �  �    C  x    D  �  �  �  +  V  �  �    8  `  �  �  	  G	  {	  �	  �	   
  `
  �
  �
  �
  7  v  �  �    P  �  �  �  .  e  �  �    H  |  �  �  )  ^  �  �    ?  v  �  �    V  �  �  �  3  m  �  <  j  �  �    :  r  �  �  "  P  �  �  	  :	  d	  �	  �	  �	  7
  q
  �
  �
    C    �  �     Y  �  �  �  4  i  �  �    J    �  �  $  Y  �  �  �  6  l  �  �    K  �  �  �  #  [  �  �  q  �  �    F  �  �  �  2  b  �  �  	  K	  {	  �	  �	  &
  ^
  �
  �
  �
  3  n  �  �    B  �  �  �    V  �  �  �  2  l  �  �    M  �  �  �  )  _  �  �    ;  r  �  �    M  �  �  �  �  �  �    H  �  �    3  \  �  �  	  K	  w	  �	  �	  +
  d
  �
  �
  �
  8  v  �  �    K  �  �  �  '  a  �  �    B  {  �  �  (  \  �  �  
  @  u  �  �     X  �  �     :  s  �  �  .  �  �  �    4  n  �  �    G  x  �  �  2	  `	  �	  �	  
  C
  u
  �
  �
    R  �  �  �  &  c  �  �    >  y  �  �  !  V  �  �    :  m  �  �    O  �  �  �  /  g  �  �    F    �  �  >  �  �  �    F  �  �    2  \  �  �  	  J	  w	  �	  �	  %
  \
  �
  �
  �
  4  p  �  �    I  �  �  �  *  a  �  �    A  y  �  �  (  _  �  �    C  y  �  �  "  [  �  �    :  s  �  �  �  �  �  �    ?  _  �  �  &  L  |  �   	  8	  i	  �	  �	  
  J
  �
  �
  �
  &  `  �  �    =  t  �  �    T  �  �  �  7  n  �  �    Q  �  �  �  1  j  �  �    L  �  �  �  .  g  �    D  �  �  �    "  P  �  �  �  5  h  �  �  	  N	  �	  �	  �	  )
  e
  �
  �
    @  {  �  �  "  W  �  �    :  p  �  �    T  �  �  �  7  o  �  �    M  �  �  �  /  h  �  �    J  �  "  g    C  �  �    7  h  �  �    X  �  �  �  /	  t	  �	  �	  
  D
  �
  �
  �
  %  `  �  �    G  �  �  �  8  m  �  �     X  �  �    >  w  �  �     [  �  �    <  v  �  �    W  �  f  �  �  B  �  �  �  #  b  �  �    H  z  �  �  	  `	  �	  �	  
  ?
  �
  �
  �
  +  f  �  �  	  C  ~  �  �  #  ^  �  �    =  v  �  �  !  W  �  �    8  m  �  �    O  �  �  �  0  i  F    �    I  _  �  �  +  ]  �  �    U  �  �  �  =	  u	  �	  �	  
  Z
  �
  �
  �
  9  q  �  �    X  �  �  �  8  r  �  �    S  �  �  �  5  n  �  �    Q  �  �  �  5  l  �  �    M  _    �  �    E  �  �  �    R  �  �    5  f  �  �  	  M	  }	  �	  �	  !
  ^
  �
  �
  �
  /  k  �  �    >  x  �  �    M  �  �  �  (  \  �  �    8  l  �  �    G  {  �  �    T  �  ]  q  �  �  �    B  z  �  �    T  �  �    1  a  �  �  	  A	  o	  �	  �	  
  O
  �
  �
  �
    W  �  �  �  #  \  �  �  �  0  g  �  �    <  r  �  �    I  }  �  �     S  �  �  �  '  �    O  �  �  �  2  m  �  �    .  b  �  �    :  h  �  �  	  G	  p	  �	  �	  
  M
  {
  �
  �
    N  �  �  �    K  �  �  �    Q  �  �  �  $  W  �  �  �  &  Z  �  �  �  (  [  �  �  �  �  9  v  �  �  �  !  p  �  �    +  \  �  �    5  W  �  �  �  /	  [	  �	  �	  �	  $
  U
  �
  �
  �
    P  �  �  �    H  |  �  �    :  t  �  �    5  h  �  �    5  c  �  �    2  �  �  B    �  �    B  m  �  �  �    L  }  �  �    8  j  �  �  �  0	  c	  �	  �	  �	  +
  ^
  �
  �
  �
  %  W  �  �  �     U  �  �  �    P  �  �  �    N    �  �    L  }  �  �    �    Y  �  �  �  �  �  "  O  u  �  �    <  n  �  �    =  f  �  �  �  7	  f	  �	  �	  �	  )
  `
  �
  �
  �
    W  �  �  �    K  �  �  �    D  y  �  �    A  s  �  �    D  q  �  �  -  S  �    I  e  �  �  �    G  |  �  �    I  u  �  �    =  l  �  �  	  3	  `	  �	  �	  �	  "
  R
  
  �
  �
    J  y  �  �    C  u  �  �    :  o  �  �    5  i  �  �     1  c  �  I  Q  -        z  �  �  �  #  D  {  �  �    6  d  �  �  �    O  �  �  �  	  D	  u	  �	  �	  
  :
  g
  �
  �
  �
  -  Z  �  �  �  &  T  �  �  �  %  X  �  �  �    T  �  �  �    N  C  �    8  d  e  |  �  �  �  �  '  q  �  �  �  �    Y  �  �  �    :  o  �  �  �  #	  X	  �	  �	  �	  
  Q
  �
  �
  �
    C  v  �  �    6  h  �  �    6  e  �  �  	  :  g  �  �      �    �  K  �  �  �  �  �      A  K  h  {  �  �  )  M  f  �  �    7  X  |  �  �  "	  K	  p	  �	  �	  	
  A
  q
  �
  �
    9  m  �  �  �  *  _  �  �  �     V  �  �  �    Q  �  �  �    2  �  f  �  �  �  �  �  �      ;  T  h  �  �  �    <  m  �  �  �    G  }  �  �  	  /	  c	  �	  �	  
  .
  Z
  �
  �
  �
  +  W  �  �  �  "  P  |  �  �    J    �  �    M  �  �  
  4  U  w  �  �  �  �  �    *  =  e  �  �  �  �    &  @  b  �  �  �  �    Y  �  �  �   	  :	  r	  �	  �	  �	  &
  a
  �
  �
  �
    S  �  �  �    L  �  �  �    E  v  �  �    H  �  �  <  t  �  �  �  �  �    '  8  d  �  �  �  �  �    3  K  h  {  �  �  �  $  H  c  �  �  	  1	  S	  u	  �	  �	  
  @
  k
  �
  �
    9  h  �  �  �  4  i  �  �  �  +  a  �  �  �  "  �  �  F  �  �  �  �  �  �         2  Y  �  �  �    7  d    �  �  �  	  ,  K  o  �  �  �  �  	  =	  |	  �	  �	  �	  -
  e
  �
  �
    ,  ]  �  �    6  c  �  �    6  e  �  �  �  2    >  r  �  �  �  �      )  D  c  �  �  �  �  
  1  W  �  �  �  �  �    ]  �  �  �  �  	  6	  j	  �	  �	  �	  
  S
  �
  �
  �
    ?  }  �  �  
  ;  s  �  �    ;  o  �  �    ?  V     [  �  �  �  �    %  =  T  l    �  �       7  X  t  �  �  �  �    5  ^  v  �  �  	  Q	  |	  �	  �	  
  I
  �
  �
  �
  	  C  �  �  �    B  }  �  �    D  z  �  �  "  M  ]  ]  ]  *  l  �  �  �  �    ,  @  S  f  w  �  �    &  @  k  �  �  �    A  i  �  �  �  	  7	  b	  �	  �	  �	   
  V
  �
  �
  �
  (  ^  �  �  �  "  Z  �  �  �  (  \  �  �  �  -  ^  �  �  �  �  C  ~  �  �  �    &  F  [  y  �  �  �    0  S  p  �  �    8  Z  �  �  �  %	  L	  v	  �	  �	  
  H
  s
  �
  �
    3  p  �  �     1  g  �  �    6  h  �  �    6  e  �  �  �  �  �  �  \  �  �  �    /  m  �  �  �  �    E  b  �  �  �    =  i  �  �  �  	  K	  z	  �	  �	  
  K
  y
  �
  �
  
  D  v  �  �    >  t  �  �  
  =  q  �  �  	  <  o  �  �    ;  G  G  G  G  �  �  �    /  U  �  �  �    7  s  �  �  �    O  |  �  �  	  5	  c	  �	  �	  �	  
  K
  ~
  �
  �
    >  }  �  �    >  v  �  �    @  s  �  �    B  s  �  �    B  t  �  �  �  �  �  �  �  �  %  Q  �  �  �  /  W  �  �  �    @  s  �  �  	  ;	  l	  �	  �	  
  3
  a
  �
  �
  �
  .  \  �  �  �    Q  �  �  �  /  a  �  �  �  0  c  �  �  �  3  i  �  �       '  '  '  '  �  �    A  t  �  �    J  s  �  �    P  �  �  �  %	  W	  �	  �	  �	  %
  V
  �
  �
  �
  $  X  �  �  �  "  W  �  �  �  !  U  �  �  �     W  �  �  �  )  ]  �  �  �  0  g  �  �  �  �  �  �    1  j  �  �    :  l  �  �    N  w  �  �  	  J	  �	  �	  �	  
  W
  �
  �
  �
  #  `  �  �  �  (  ]  �  �    3  g  �  �    6  i  �  �    8  t  �  �    A  v  �  �    8  W  g  �    L  �  �  �  *  X  �  �    @  m  �  �  	  J	  |	  �	  �	  
  P
  �
  �
  �
  %  Z  �  �    7  l  �  �    E  �  �  �    T  �  �  �  "  X  �  �  �  2  h  �  �    6  k  �  �    �  �    W  �  �  �    L  �  �    0  ]  �  �  	  N	  z	  �	  �	  +
  e
  �
  �
     >  |  �  �    V  �  �  �  4  r  �  �    Q  �  �  �  4  i  �  �    H  }  �  �  $  [  �  �    <  �  �  �  3  }  �  �    >  s  �  �  2  ^  �  �  	  H	  y	  �	  �	  '
  e
  �
  �
    B  �  �  �    [  �  �    :  u  �  �  "  W  �  �  	  ?  s  �  �  #  [  �  �    =  u  �  �    V  �  �  �    7  �  �    ,  W  �  �    E  t  �  �  -	  _	  �	  �	  �	  ?
  v
  �
  �
    Q  �  �  �  (  d  �  �    @  y  �  �  $  X  �  �    =  q  �  �    V  �  �  �  4  n  �  �    .  �  �    6  u  �  �  )  ]  �  �    @  p  �  �   	  W	  �	  �	  �	  3
  n
  �
  �
    K  �  �  �  +  d  �  �    D  �  �  �  .  d  �  �    L  �  �  �  ,  f  �  �    H  �  �  �  ,  m  �  �    O  �  �  �     G  �  �    <  e  �  �  	  W	  �	  �	  �	  1
  m
  �
  �
    I  �  �  �  '  a  �  �    C  |  �  �  *  `  �  �    F  |  �  �  )  b  �  �  
  E  ~  �  �  &  �  h  �  �  !  i  �  �    7  g  �  �     S  �  �  �  6	  n	  �	  �	  
  O
  �
  �
  �
  -  f  �  �    E  ~  �  �  &  ^  �  �  
  A  y  �  �  "  Z  �  �    <  u  �  �    W  �  �  �  ^  �  �  �    3  l  �  �  +  [  �  �    L  �  �  �  .	  e	  �	  �	  
  I
  �
  �
  �
  +  e  �  �    K  �  �  �  *  c  �  �    I  �  �  �  0  h  �  �    L  �  �  �  /  h  �  �    P  )  &    7  g  �  �  �  9  Y  �  �    R  |  �  �  8	  q	  �	  �	  
  R
  �
  �
  �
  .  l  �  �    I  �  �  �  (  b  �  �    F  ~  �  �  .  d  �  �    J  �  �  �  +  e  �  �    b  �      S  ;  �  �  �  0  Q  �  �    L  �  �  �  9	  n	  �	  �	  
  G
  
  �
  �
    X  �  �  �  /  k  �  �    D  �  �  �  &  ]  �  �  
  >  s  �  �  "  X  �  �    ;  r  �  �  �  �  z  �       X  �  �  �  C  �  �  �  )  ]  �  �  	  :	  g	  �	  �	  
  L
  |
  �
  �
  *  i  �  �    H  �  �  �  &  f  �  �    I  �  �  �  2  i  �  �    S  �  �    <  s  �  �  �  �  O  �  �  �  2  �  �  �    >  �  �  �    O  �  �  	  H	  z	  �	  
  B
  q
  �
  �
  ,  k  �  �    O  �  �  �  0  n  �  �    R  �  �    ;  v  �  �  !  [  �  �    ;  u  �  �  B    <  r  �  �  �  ,  g  �  �    D  �  �  	  7  o  �  �  +	  Z	  �	  �	  
  K
  |
  �
  �
  /  k  �  �    O  �  �  �  ,  j  �  �    J  �  �  �  0  h  �  �    O  �  �  �  6  n  �  Z  �  �  <  k  �  �  �  8  p  �  �    C  |  �  �  &  X  �  �  �  0	  e	  �	  �	  

  @
  v
  �
  �
    N  �  �  �  %  [  �  �     4  i  �  �    C  x  �  �    R  �  �  �  )  `  �  �  �  �  �  �  "  p  �  �  �    ]  �  �    ,  `  �  �    D  l  �  �  *	  Y	  �	  �	  �	  ,
  f
  �
  �
  �
  -  j  �  �    7  s  �  �    D  {  �  �     R  �  �  �  +  ^  �  �  �  3  h  B  h  �  �  �  *  �  �  �  �  1  h  �  �    4  m  �  �  $  J  m  �  �  *	  X	  	  �	  �	  "
  b
  �
  �
  �
  !  ^  �  �  �  "  ^  �  �     .  a  �  �    5  d  �  �    >  l  �  �      N  �  �  �    '  �  �  �  �  @  d  �  �    4  q  �  �    B  f  �  �  	  G	  q	  �	  �	  
  E
  u
  �
  �
  �
  3  s  �  �  �  .  c  �  �  �  '  ^  �  �  �  ,  W  �  �  �  -  [  �  �  O  �  �  �    =  �  �  �    B  ~  �  �    =  l  �  �    A  k  �  �  	  :	  l	  �	  �	  
  6
  e
  �
  �
  �
  -  c  �  �  �  (  ]  �  �  �  #  W  �  �  �  !  R  �  �  �    N  �  �  B  �  �  �    9  u  �  �  �    M  �  �  �    D  {  �  �    ;  j  �  �  	  0	  a	  �	  �	  �	  +
  [
  �
  �
  �
  "  R  �  �  �    Q  �  �  �    M  ~  �  �    I  {  �  �    =  '  _  �  �  �  �  �  E  �  �  �    ,  [  �  �  �    =  s  �  �  �  /  g  �  �  �   	  R	  �	  �	  �	  
  F
  |
  �
  �
  
  :  p  �  �    6  g  �  �  	  8  e  �  �    7  e  �  �  �  G  s  �  q  �  �  �  L  l  `  �  �  �    A  X  �  �  �  /  U    �  �    R  ~  �  �  	  E	  v	  �	  �	  �	  1
  e
  �
  �
  �
  #  Y  �  �  �    M  �  �  �    K  �  �  �    G  z  �  c  h  �  �  �    �    �  ,  /  i  �  �      I    �  �    2  c  �  �     %  P  �  �  �  $	  P	  ~	  �	  �	  
  J
  u
  �
  �
    =  i  �  �  �  2  d  �  �  �  1  j  �  �  �  +  c  w  ~  �  �  �  �  �  �  �  -    e  �  �  �  �    _  �  �  �  �  *  d  �  �  �    E  �  �  �  �  ,	  f	  �	  �	  �	  *
  ^
  �
  �
  �
  $  S  �  �  �  !  K  {  �  �    O  {  �  �    {  �  �  �  �  �  �  �  �  :  _  z  �  �  �  �    =  Z  z  �  �  �  .  Z  x  �  �    D  j  �  �  �  1	  a	  �	  �	  �	  
  X
  �
  �
  �
    K  �  �  �    ;  r  �  �    9  p  �  �  w  �  �  �  �  �  �    $  I    �  �  �  �  �    $  /  M  q  �  �    %  C  }  �  �    3  [  �  �  �  "	  K	  |	  �	  �	  #
  J
  v
  �
  �
     M  v  �  �    L  z  �  �  
  D  {  �  �  �  �  �  �  �  �  �    I  �  �  �  �       =  ^  ~  �  �  �       P  z  �  �  �  �  
  J  �  �  �  �  2	  o	  �	  �	  �	  &
  d
  �
  �
    /  b  �  �    1  _  �  �    4  `  �  �  �  �  �  �  �    (  ^  �  �  �  �    /  X  s  �  �  �  �  '  E  c  ~  �  �  �    /  Z  x  �  �  �  1	  e	  �	  �	  �	  #
  c
  �
  �
  �
    Y  �  �  �    V  �  �  �  %  S  �  �  �  �  �        1  I  �  �  �  �  	  &  ?  T  h  z  �  �  �     7  Q  �  �    F  b  �  �  �  	  O	  	  �	  �	  

  C
  w
  �
  �
  �
  1  l  �  �  �  /  f  �  �     1  b  �  �    
  �          )  ;  V  �  �  �    %  c  �  �  �  �    2  U  z  �  �    +  B  c  �  �  	  H	  p	  �	  �	  
  H
  |
  �
  �
    F  �  �  �    E  �  �  �    J  �  �  �  '  6  6  6    +  5  <  M  _  �  �  �  �    1  [  �  �  �    ;  v  �  �  	  .  ]  �  �  �  �  '	  Z	  �	  �	  �	  
  F
  �
  �
  �
    L  |  �  �    I    �  �    N  �  �  �    O  �  �  �  �  4  d  x  �  �  �  �      A  e  �  �  �  $  M  n  �  �    ;  b  �  �  �  '	  N	  x	  �	  �	  
  A
  l
  �
  �
    ,  h  �  �    1  i  �  �    2  f  �  �    @  p  �  �  �  �  �  �  N  �  �  �      7  Q  h  �  �    0  T  ~  �  �    ?  q  �  �  �  ,	  `	  �	  �	  �	  "
  W
  �
  �
  �
    T  �  �  �    M  �  �  �    G  |  �  �    B  w  �  �    J  a  a  a  a  �  �  �    1  [  v  �  �  �  !  G  n  �  �    :  j  �  �  �  3	  e	  �	  �	  �	  (
  `
  �
  �
  �
  )  ]  �  �  �  (  Y  �  �  �  (  W  �  �  �  &  U  �  �  �  #  S  �  �  �  �  �  �  �  �  �    F  �  �  �  #  M  n  �  �  �    T    �  �  	  U	  �	  �	  �	  +
  b
  �
  �
  �
  8  o  �  �    ;  q  �  �    G  }  �  �    K  �  �  �    N  �  �  �    R  �  �  �  �  �  �  �    Q  �  �    3  f  �  �    8  q  �  �  �  *	  b	  �	  �	  �	  +
  g
  �
  �
    9  p  �  �    E  }  �  �    P  �  �  �  (  ]  �  �    7  k  �  �    G  ~  �  �    -  /  �  �      h  �  �    >  p  �  �  4  W  �  �  �  1	  e	  �	  �	  
  5
  d
  �
  �
    :  l  �  �  	  ;  p  �  �    K  ~  �  �    S  �  �  �  (  b  �  �     5  k  �  �    A  x  �  �  �    e  �  �  �  !  X  �  �     3  g  �  �  	  C	  u	  �	  �	  
  P
  �
  �
  �
  !  ^  �  �  �  0  i  �  �    A  y  �  �    L  �  �  �     T  �  �  �  1  e  �  �    :  n  �  �  �  �  �    U  �  �    -  g  �  �    J  �  �  	  :	  h	  �	  �	  
  L
  �
  �
  �
  !  ^  �  �  �  1  n  �  �    H  �  �  �  $  _  �  �    9  s  �  �    K  �  �  �  )  `  �  �    �  �  �    V  �  �    *  b  �  �    J  |  �  �  9	  f	  �	  �	  
  L
  �
  �
  �
  "  b  �  �    =  {  �  �    W  �  �    :  q  �  �     U  �  �    :  o  �  �    S  �  �  �  1  �  �  �  �  4  ~  �  �     L  �  �    ;  f  �  �  	  P	  �	  �	  �	  0
  i
  �
  �
    D    �  �    X  �  �  �  3  m  �  �    K  �  �  �  /  d  �  �    G  }  �  �  '  _  �  �    �  �  �    5  s  �  �    ?  �  �    5  c  �  �  	  N	  ~	  �	  �	  +
  e
  �
  �
    ?  y  �  �    W  �  �  �  5  p  �  �    U  �  �    9  o  �  �    R  �  �  �  2  k  �  �      �  �  	    }  �  �    =  �  �    1  [  �  �  	  M	  |	  �	  �	  *
  e
  �
  �
    B  }  �  �    [  �  �    :  u  �  �     V  �  �    <  r  �  �    W  �  �  �  9  r  �  �      �  �  �    U  �  �    .  a  �  �    I  }  �  �  +	  c	  �	  �	  
  ?
  z
  �
  �
    S  �  �  �  5  k  �  �    O  �  �  �  4  k  �  �    K  �  �  �  ,  f  �  �    F  �  �  �  �  5  �  �    -  h  �  �  !  R  �  �  �  @  r  �  �  	  Q	  �	  �	  �	  &
  j
  �
  �
    F  �  �    6  l  �  �     X  �  �    ?  w  �  �  #  ]  �  �    A  z  �  �  $  ]  �  �    �  �  �  �  �  7  �  w  �  &  H  z  �  �  '  Z  �  �  �  E	  �	  �	  �	  )
  n
  �
  �
    M  �  �  �  .  k  �  �    M  �  �  �  ,  e  �  �    C  z  �  �  %  \  �  �    ?  v  �  �  �  B  �  �  �  #  .  Z  �  �    V  �  �    P  z  �  �  0	  i	  �	  �	  
  E
  x
  �
  �
  %  _  �  �    A  |  �  �  "  \  �  �    >  x  �  �    P  �  �  �  0  h  �  �    J  �  �    Q    8  �  �  �  :  e  �  �  .  `  �  �    B  }  �  �  /	  g	  �	  �	  
  >
  {
  �
  �
  #  \  �  �    E  }  �  �  /  i  �  �    R  �  �  �  :  s  �  �  "  \  �  �  	  D    �  >  k  �  .  �  �  �    T  �  �  �  )  h  �  �    V  �  �  	  ?	  z	  �	  �	  2
  p
  �
  �
    [  �  �  	  @  {  �  �  +  c  �  �    R  �  �    <  r  �  �    S  �  �  �  ;  v  �  �  �  �  �  =  U  �  �    N  �  �    =  z  �  �  (  c  �  �  	  J	  �	  �	  �	  1
  k
  �
  �
    U  �  �    ;  r  �  �     Y  �  �    >  v  �  �    F  {  �  �    R  �  �  �  '  �  �  �  �  �  ;  l  �  �    A  |  �  �    N  �  �  �  0  b  �  �  	  A	  s	  �	  �	  
  N
  �
  �
  �
    Z  �  �  �  -  f  �  �  
  <  s  �  �    K  �  �  �  '  Z  �  �  �  3  h  /  S  s  �  �  �  3  b  �  �  �  /  p  �  �  
  7  s  �  �    G  w  �  �  +	  Y	  �	  �	  �	  5
  g
  �
  �
  �
  8  r  �  �  	  A  {  �  �    K  �  �  �    T  �  �  �  )  ]  �  �  �  �    7  q  �  �     L  �  �  �  �  ;  �  �  �    :  z  �  �     I  t  �  �  &	  S	  }	  �	  �	  )
  Y
  �
  �
  �
  $  X  �  �  �  )  ^  �  �  �  -  _  �  �  �  /  `  �  �  �  /  `  �  �  �    \  �  �  �  �  J  �  �  �  �  3  w  �  �    &  _  �  �    0  Q  �  �  �  )	  X	  ~	  �	  �	  #
  T
  �
  �
  �
    N    �  �    E  y  �  �    <  q  �  �    4  i  �  �    �  �    F  �  �  �    ?  n  �  �  �    N  w  �  �    <  i  �  �     4  d  �  �  �  -	  a	  �	  �	  �	  #
  Y
  �
  �
  �
    S  �  �  �    M  �  �  �    I  |  �  �    I  x  �  �  �  �    k  d  �  �  �  �    :  q  �  �    2  k  �  �    9  _  �  �    7  [  �  �  �  .	  ^	  �	  �	  �	  "
  Y
  �
  �
  �
    O  �  �  �    A  ~  �  �    :  q  �  �    :  i  �  �    =  �  %  9  P  �  �  �    <  �  �  �    4  j  �  �    7  c  �  �    /  Y  �  �  �  	  K	  x	  �	  �	  
  F
  r
  �
  �
    @  o  �  �     8  m  �  �  �  /  g  �  �  �  '  ]  �  !    �  �  �  *  n  �  �  �    8  {  �  �  �  '  ^  �  �  �    F    �  �    7  m  �  �   	  *	  Z	  �	  �	  �	  
  K
  
  �
  �
    D  r  �  �    K  v  �  �    K  x  �  �      �  �  �    �  3  f    �  �  �  )  \  z  �  �  �    L  q  �  �  �  .  _  �  �  �    L  �  �  �  
	  D	  {	  �	  �	  �	  1
  i
  �
  �
  �
  "  X  �  �  �     R  �  �  �  &  Q  �  �  �  �  �  �  �  3  I  U  �  �  �  �    #  1  S  h  �  �    .  F  z  �  �    :  f  �  �    /  T  �  �  �  1	  Y	  �	  �	  �	  +
  Y
  �
  �
  �
    O  �  �  �    H  ~  �  �    @  |  �  �  �  �  �  C  `  �  �  �  �  �  �  �  �    <  �  �  �  �    V  �  �  �  �  *  e  �  �  �    H  �  �  �  	  >	  w	  �	  �	  
  ?
  p
  �
  �
    <  e  �  �    B  l  �  �    E  �  �  �  �  %  T  q  �  �  �  �  �       C  o  �  �  �  �    9  a  {  �  �  �  �  @  l  �  �  �  %  ^  �  �  �  	  [	  �	  �	  �	  
  R
  �
  �
  �
    K  �  �  �    E  }  �  �  &  �  �  �    V  s  �  �  �  �      ;  P  ]  �  �  �       ?  U  m  �  �  �  �    <  H  w  �    :  [  }  �  �  8	  k	  �	  �	  �	  0
  o
  �
  �
  �
  ,  k  �  �  �  *  f  �  �  	  3    �  �  7  m  �  �  �  �  �      )  4  L  �  �  �      _  �  �    '  Q  v  �  �  �    K  `    �  �  2	  ^	  �	  �	  �	  ,
  [
  �
  �
  �
    [  �  �  �    Y  �  �  �  #  V  �  b  ]  c    �  �  �  �  8  ^  x  �  �  �  �    #  H  f  �  �  �    +  ]  �  �    A  d  �  �  	  D	  w	  �	  �	  �	  4
  f
  �
  �
  �
    T  �  �  �     S  �  �  �  #  M  �  �  �  �  �  �  �  �  �  �    .  r  �  �  �    B  r  �  �  �    .  T  {  �  �    +  G  m  �  �  	  B	  n	  �	  �	  
  <
  p
  �
  �
     ;  r  �  �    ;  v  �  �    C  z  �  �    .  .  .  �  �  �  �      R  �  �  �    9  g  �  �  �    M  �  �  �    =  l  �  �  �  	  I	  z	  �	  �	   
  4
  h
  �
  �
  �
  8  m  �  �    5  k  �  �    :  n  �  �    8  k  �  �  �  �  �  �  �  
  @  x  �  �  �     A  s  �  �    H  r  �  �    A  j  �  �  	  7	  e	  �	  �	  
  0
  _
  �
  �
  �
    M  �  �  �    M  �  �  �     Q  �  �  �  $  _  �  �  �    (  (  (  �  �    N  ~  �  �    %  \  �  �     -  V  �  �  �  %  [  �  �  �  '	  \	  �	  �	  �	  )
  ]
  �
  �
  �
  #  ^  �  �  �  %  \  �  �  �  %  [  �  �  �  %  Z  �  �  �  (  c  �  �  �  �      P  �  �  �    5  j  �  �    ;  f  �  �    A  m  �  �  	  =	  o	  �	  �	  
  >
  v
  �
  �
    A  y  �  �    D  {  �  �    I  }  �  �    M  �  �  �    P  �  �  �     R  �  1  w  �  �  �    %  W  �  �    4  g  �  �     L  z  �  �  ,	  ^	  �	  �	  �	  6
  m
  �
  �
    A  z  �  �    N  �  �  �  %  \  �  �  �  +  a  �  �  �  1  g  �  �    7  l  �  �    F  �  �  �    3  e  �  �    +  L  x  �    7  j  �  �  	  W	  �	  �	  �	  7
  s
  �
  �
    P  �  �  �  -  i  �  �    F  �  �  �  +  `  �  �    E  z  �  �  %  ]  �  �    <  u  �  Z  �  �  �     _  �  �    -  b  �  �    6  f  �  �  	  <	  m	  �	  �	  

  F
  }
  �
  �
    X  �  �  �  -  l  �  �    E  ~  �  �  '  \  �  �    ?  t  �  �    V  �  �  �  5  n  �  �  �  �    G  �  �  �  #  S  �  �    8  b  �  �  	  C	  s	  �	  �	  
  J
  {
  �
  �
    Y  �  �  �  )  `  �  �  	  ?  u  �  �    J  ~  �  �  !  V  �  �  �  6  l  �  �    C  y  �  �  �    o  �  �  �    Y  �  �    7  i  �  �  /  \  �  �  	  @	  u	  �	  �	  
  V
  �
  �
  �
  3  o  �  �    O  �  �  �  4  n  �  �    R  �  �  �  5  o  �  �    R  �  �  �  8  q  �  �  �  G  �  �  �    L  �  �    9  n  �  �  )  Z  �  �  
	  F	  y	  �	  �	  $
  `
  �
  �
     <  y  �  �    V  �  �    8  q  �  �    T  �  �    ;  q  �  �    W  �  �  �  9  r  �  �  �    V  �  �    E  }  �  �  3  c  �  �    N  �  �  �  .	  h	  �	  �	  
  H
  �
  �
  �
  &  `  �  �    @  y  �  �  "  Z  �  �    =  t  �  �    X  �  �    :  s  �  �    U  h  �    f  �  �  �    N  �  �    D  |  �  �  ,  _  �  �  	  F	  z	  �	  �	  +
  b
  �
  �
    I  �  �  �  &  `  �  �    F  �  �  �  -  e  �  �    K  �  �  �  .  f  �  �    J  �  x  /  :  q  z  �       i  �  �    C  u  �    <  k  �  �  	  T	  �	  �	  �	  4
  n
  �
  �
    L  �  �  �  (  f  �  �    D    �  �  +  a  �  �    H  ~  �  �  ,  c  �  �    G  �  �  p  �  >  �  �  �    e  �  �    X  �  �    8  h  �  �  	  G	  y	  �	  �	  
  X
  �
  �
  �
  0  j  �  �  	  D  �  �  �  !  [  �  �    7  p  �  �    Q  �  �  �  6  l  �  �    P  Q    �  0  �  �  �    i  �  �  �  ,  f  �  �  	  4  g  �  �  	  H	  w	  �	  �	  2
  e
  �
  �
    P  �  �  �  -  n  �  �    M  �  �  �  1  l  �  �    S  �  �    <  s  �  �  !  Z  J  �  �  �  U  �  �  �    `  �  �  �    L  �  �    =  t  �  	  6	  g	  �	  �	  1
  b
  �
  �
    Q  �  �  �  1  o  �  �    R  �  �     ;  v  �  �  "  \  �  �    <  v  �  �    V  R  �  �  �  K  �  �  �  �    >  �  �    :  �  �  �  /  r  �  �  /	  b	  �	  �	  
  D
  {
  �
  �
  (  `  �  �    I  �  �  �  ,  d  �  �    F  t  �  �    S  �  �  �  7  p  �  �    _  �  ^  v  �  �  4  �  �  �  &  �  �  �    X  �  �    9  l  �  �  	  F	  y	  �	  �	  )
  d
  �
  �
    J  �  �  �  -  n  �  �    Y  �  �    F  �  �  �  8  r  �  �  *  f  �  �    }  �  I  }  �  �    n  �  �  �  9  z  �  �    E  �  �  	  =  r  �  �  =	  s	  �	  �	  '
  f
  �
  �
    N  �  �  �  6  t  �  �     [  �  �    F  �  �  �  5  l  �  �  "  \  �  �    �  �  (  ^  �  �  �    W  �  �  �  2  �  �  �  )  `  �  �    L  �  �  �  9	  m	  �	  �	   
  \
  �
  �
    C  }  �  �  "  `  �  �    A  ~  �  �  )  a  �  �    J  �  �  �  2  k  �  �  �  �    T  }  �  �    V  �  �  �    [  �  �    3  i  �  �    >  x  �  �  	  O	  �	  �	  �	  +
  _
  �
  �
    8  m  �  �    E  z  �  �    R  �  �  �  *  `  �  �    7  m  �    �  �  �    ^  }  �  �  �  2  y  �  �  �  6  y  �  �    @  {  �  �  +  T  �  �  �  8	  f	  �	  �	  
  <
  r
  �
  �
    F    �  �    O  �  �  �  %  Y  �  �  �  1  d  �  �    :  '  L  �  �  �  �  N  �  �  �  
  ?  �  �  �    E  {  �  �    A  ~  �  �  *  Q  |  �  �  3	  a	  �	  �	  �	  0
  j
  �
  �
  �
  2  l  �  �    4  l  �  �    7  k  �  �    ?  o  �  �    ,  f  �  �  �    T  �  �  �  	  3    �  �    3  f  �  �    2  b  �  �    B  b  �  �  	  F	  p	  �	  �	  �	  >
  t
  �
  �
  �
  -  m  �  �  �  "  ]  �  �  �    R  �  �  �  '  N  �     H  }  �  �  �  <  �  �  �  �  7  ~  �  �    *  m  �  �    2  _  �  �  
  9  _  �  �  	  3	  _	  �	  �	  �	  0
  a
  �
  �
  �
  (  ]  �  �  �     V  �  �  �    M  �  �  �    I  y  �  ;  �  �  �  �  9  t  �  �  �    \  �  �  �    G  �  �  �    2  k  �  �  �  &  Y  �  �  �  "	  Q	  �	  �	  �	  
  F
  x
  �
  �
    E  t  �  �    D  p  �  �    A  m  �  �  �  d  �  2  s  �  �  �  �  J  v  �  �  �  )  W  |  �  �    ;  g  �  �  �  *  _  �  �  �    J  ~  �  �  �  :	  s	  �	  �	  �	  '
  d
  �
  �
  �
    U  �  �  �  #  N  �  �  �  &  O  }  �  �    B  2  M  �  �  �  5  ;  T  m  �  �    )  G  p  �  �    6  d  �  �    9  b  �  �    7  ]  �  �  �  #	  T	  z	  �	  �	  
  J
  z
  �
  �
    B  |  �  �  �  7  s  �  �     .  f    /  K  g  {  �  �  �  �  �      Z  �  �  �  �  -  o  �  �  �    K  �  �  �    2  h  �  �  
  0  `  �  �  	  .	  X	  �	  �	  �	  (
  O
  |
  �
  �
  $  U  }  �  �  $  Z  �  �  �    A  l  H  M  �  �  �  �  �  �  �  �  C  l  �  �  �    Q  �  �  �  �    L  ~  �  �  �  0  l  �  �  �    [  �  �  �  	  N	  �	  �	  �	  
  @
  |
  �
  �
    7  m  �  �    ?  l  �  �  m  �  x  �  �  �  �  �  �  �    F  b  y  �  �  �    ;  N  ^  m  �  �    :  Q  x  �  �  0  O  o  �  �  /  c  �  �  �  %	  d	  �	  �	  �	  
  \
  �
  �
  �
    R  �  �  �    O  �  �  �  �  �  �  �  �  �  �  �    $  u  �  �  �  �      ,  @  Q  f  �  �  �  
  *  r  �  �  $  ;  h  �  �  1  S  u  �  �  4	  h	  �	  �	  �	  /
  n
  �
  �
  �
  *  l  �  �  �  )  h  �  �  �  �  �  �  �  �  �  �      :  t  �  �  �    `  �  �  �  �    1  H  s  �  �      "  L  �  �    7  W  �  �  	  >	  i	  �	  �	  �	  ?
  r
  �
  �
  �
  ;  y  �  �    <  z  �  �    �  �  �  (  G  P  \  l  �  �  �  �  �    .  i  �  �  �    >  �  �      A  w  �  �  �    J  t  �  �  �  /	  ]	  �	  �	  �	  %
  N
  �
  �
  �
    O  �  �  �    O  �  �  �    L  �  �  ,  O  z  �  �  �  �      ,  ?  o  �  �    &  S  ~  �  �  �    A  o  �  �    F  m  �  �   	  Q	  y	  �	  �	  
  X
  �
  �
  �
    9  p  �  �    <  o  �  �    C  d  �  �  �  �  �  B  �  �  �  �    8  J  f  �  �  �    2  V  �  �  �  *  T  �  �  �    D  n  �  �  	  8	  q	  �	  �	  �	  1
  h
  �
  �
  �
  ,  f  �  �  �  0  e  �  �  
  :  l  �  �    F  U  U  U  B  y  �  �  �  �  C  �  �  �    -  Q  m  �  �  �  (  O    �  �  ,  ^  �  �  �  .	  a	  �	  �	  �	  -
  [
  �
  �
  �
  +  c  �  �    5  g  �  �    7  x  �  �    P  �  �  �           `  �  �  �  �  <  �  �  �    1  n  �  �    ;  c  �  �  �    O  ~  �  �  	  N	  �	  �	  �	  !
  Y
  �
  �
  �
  &  _  �  �  �  4  k  �  �  
  @  v  �  �    K  �  �  �  &  _  �  �  �  k  �  �    g  \  �  �      X  �  �    3  c  �  �    ?  q  �  �  	  6	  p	  �	  �	  
  4
  k
  �
  �
    ;  t  �  �    C  {  �  �    N  �  �  �  &  Y  �  �  �  2  j  �  �    C  �  �  �  (  }  �  �  �  (  y  �  �  �  -  e  �  �    <  l  �  �  	  C	  u	  �	  �	  
  K
  ~
  �
  �
    Q  �  �  �     U  �  �  �  '  \  �  �  �  /  c  �  �    7  k  �  �  	  ?  v  �  �  �  %  v  �  �  �  %  s  �  �    ;  y  �  �  (  S  �  �  		  =	  j	  �	  �	  
  N
  
  �
  �
    \  �  �  �  .  j  �  �  	  ?  s  �  �    I  ~  �  �     T  �  �  �  *  ^  �  �  �  �  �    \  �  �    5  f  �  �  %  P  �  �    @  l  �  �  &	  ]	  �	  �	  
  B
  |
  �
  �
    ]  �  �    ;  y  �  �  "  Z  �  �  
  A  x  �  �  %  ]  �  �    @  x  �  �  !  [  �  �    �  G  �  �  	  -  g  �  �    L  �  �    E  z  �  �  :	  l	  �	  �	  
  [
  �
  �
  �
  ;  x  �  �    Z  �  �    <  w  �  �  $  Z  �  �    D  z  �  �  +  b  �  �    G  w  �  �     u  �  �  �    X  �  �  �  ,  d  �  �    =  p  �  �  	  V	  �	  �	  �	  7
  p
  �
  �
    N  �  �  �  +  h  �  �    F  �  �  �  (  _  �  �    B  x  �  �  "  [  �  �    4  �  �    j  �  �  �    U  �  �    .  d  �  �  %  R  �  �  �  8	  l	  �	  �	  
  N
  �
  �
  �
  ,  g  �  �  
  D  �  �  �  &  _  �  �    B  z  �  �  '  \  �  �    ?  v  �  �  $  \  �  �  �  C  �  �  �    I  �  �    /  i  �  �    P  �  �  	  =	  o	  �	  �	  
  X
  �
  �
  �
  6  q  �  �    P  �  �  �  0  j  �  �    L  �  �  �  2  h  �  �    M  �  �  �  .  h  �  �  �    S  �  �    >  x  �  �  )  [  �  �    C  w  �  �  	  Z	  �	  �	  �	  0
  p
  �
  �
    G  �  �  �  +  a  �  �    H  }  �  �  .  e  �  �    I  �  �  �  (  c  �  �  
  C  �  �    `  z  �  �    I  _  �    4  i  �  �    K  �  �  �  '	  i	  �	  �	  
  G
  �
  �
  �
  .  k  �  �    T  �  �    =  u  �  �  #  \  �  �    A  y  �  �  %  ^  �  �    A  z        m    h  �  	  G  b  �  �    U  �  �    J  �  �  �  4	  x	  �	  �	  
  \
  �
  �
    @  z  �  �    [  �  �    :  u  �  �    T  �  �     6  m  �  �    P  �  �  �  3  j  �  �  �  )  +  f  �  �    Z  �  �    X  �  �  �  A  �  �  �  #	  [	  �	  �	  �	  4
  i
  �
  �
    C  y  �  �  #  Z  �  �     :  r  �  �    K  �  �  �  )  c  �  �    C  |  �  �  %  �  �  �  �  G  +  k  �    L  o  �  �  3  a  �  �  �  ;  u  �  �  	  D	  �	  �	  �	  $
  `
  �
  �
    E  �  �  �  1  k  �  �    S  �  �    ;  t  �  �  $  ]  �  �    G  �  �  �  /  �  �  �  �  �  /  o  �  �    M  l  �  �    J  �  �    B  w  �  �  6	  u	  �	  �	  
  Z
  �
  �
    =  z  �  �  &  a  �  �    P  �  �    ?  z  �  �  ,  g  �  �    M  �  �  �  1  �    d  �  �  *  '  E  �  �     B  �  �    =  o  �  �  "  b  �  �  	  Q	  �	  �	  
  @
  z
  �
  �
  "  `  �  �  	  E    �  �  -  h  �  �    U  �  �    F  �  �  �  7  r  �  �    �  3  	  -  �  �  �  0  p  �  �    Z  �  �    M  �  �  	  ?  t  �  �  8	  p	  �	  �	  .
  l
  �
  �
    P  �  �  �  2  t  �  �  %  _  �  �    O  �  �    B  {  �  �  3  o  �  �  #    8  �    O  �  �  �  1  b  �  �    _  �  �     ]  �  �    Y  �  �  	  Q	  �	  �	  
  G
  �
  �
  �
  9  y  �  �  '  g  �  �    P  �  �    ;  y  �  �  -  e  �  �    U  }  �  �  �  �  �  �  -  ?  �  �  �  3  s  �  �  &  _  �  �    P  �  �    ?  u  �  �  '	  _	  �	  �	  

  C
  �
  �
  �
  0  f  �  �    C  w  �  �    P  �  �  �    T  �  �  �  )  `  �  �  �  �  �  w  �  �    K  �  �  �  *  _  �  �     5  m  �  �    G  |  �  �  #  W  �  �  �  .	  f	  �	  �	  �	  8
  s
  �
  �
    C  ~  �  �    O  �  �  �  *  ]  �  �    8  k  �  �    E  �    N  y  �  �    @  |  �  �    F  �  �  �    H  �  �  �     L  �  �    3  ]  �  �  	  ?	  l	  �	  �	  
  H
  |
  �
  �
    Q  �  �  �    X  �  �  �  (  _  �  �  �  0  e  �  �  �  �    ]  z  �  �    Y  �  �  �    S  �  �  �    O  �  �  �    G  �  �  �  )  O  �  �  �  -	  Y	  �	  �	  �	  *
  Y
  �
  �
  �
  /  a  �  �  �  /  b  �  �  �  /  `  �  �  �  .  ^    �  �    b  �  �  �    U  �  �  �    H  �  �  �  �  2  p  �  �       Y  �  �  �  &  L  �  �  �  $	  O	  x	  �	  �	  
  M
  y
  �
  �
    C  v  �  �    ;  m  �  �  �  3  e  �  �  X  z  �  %  s  �  �  �    C  j  �  �  �    H  r  �  �    1  `  �  �  �  +  T  �  �  �  "  U  ~  �  �  	  M	  �	  �	  �	  

  E
  ~
  �
  �
    9  u  �  �    1  h  �  �    1  `  �  Y  i  �    X  \  t  �  �  �    1  d  �  �  �    U  �  �  �    F  |  �  �  "  ;  h  �  �    G  _  �  �  	  J	  r	  �	  �	  
  A
  v
  �
  �
  �
  0  n  �  �  �     `  �  �  �    P  ^  �  �  �  �      F  �  �  �  �  %  m  �  �  �    O  �  �  �    E  �  �  �    ?  m  �  �  
  0  ]  �  �  	  /	  V	  �	  �	  �	  -
  V
  }
  �
  �
  (  Z  �  �  �    U  �  �  �    �  �  �  e  z  �  �    P  �  �  �  �  (  r  �  �  �    J  �  �  �  �  +  m  �  �  �    X  �  �  �    @  |  �  �   	  .	  i	  �	  �	   
  &
  X
  �
  �
  	  0  Z  �  �  	  9  _  �  �    �  �  �  �  �  |    /  l  t  �  �    I  _  r  �  �  �  1  O  l  �  �    D  `  �  �     E  n  �  �  �  :  s  �  �  �  ,	  j	  �	  �	  �	  
  ^
  �
  �
  �
    V  �  �  �  #  S  �  :    �  s  �  �    *  :  [  w  �  �        3  3  �  �  �      [  �  �  	    L  �  �    4  X  �  �    L  e  �  �  	  N	  {	  �	  �	  
  G
  �
  �
  �
  �
  >  �  �  �    <  |  V  =  �  �  �  �  &  O  �  �  �  �  �  �  �    
  ,  o  �  �  �  �  P  �  �  �    D  �  �    )  L  �  �    B  c  �  �  	  P	  y	  �	  �	  
  T
  �
  �
  �
    R  �  �  �    P  �  i  O  ?  2  0  9  ^  �  �  �  �  &  6  U  l  �  �  �  �    2  L  �  �  �  �  	  G  �  �      E  �  �    7  W  �  �  	  F	  o	  �	  �	  	
  L
  �
  �
  �
    J  �  �  �    K  �  �  �  }  w  z  �  �  �  �  �    (  g  �  �  �  �  L  {  �  �  �    5  W  |  �  �    )  5  a  �  �    ;  ^  �  �  	  9	  f	  �	  �	  �	  9
  j
  �
  �
  �
  5  r  �  �    8  t  �  �    �  �  �  �  �  �  �  %  _  �  �  �  �    R  �  �  �  �  #  \  �  �  
  +  T  �  �  �    A  u  �  �  �  )	  `	  �	  �	  �	  
  W
  {
  �
  �
    @  y  �  �    B  y  �  �    =  q  �  �  �  �  �  �    E  v  �  �  �    \  �  �    )  ]  �  �  �  #  Q  �  �  �    S  �  �  �  #	  Z	  �	  �	  �	  
  T
  �
  �
  �
  $  ^  �  �    ,  _  �  �    ;  k  �  �  �        �  �  "  S  f  �  �  �  �    A  �  �  �    F  �  �  �  -  [  �  �    F  t  �  �  	  I	  �	  �	  �	  $
  \
  �
  �
    :  m  �  �    F  {  �  �    W  �  �  �  &  Z  �  �  �  �  �    %  L  �  �  �  �  �    I  �  �  �    M  �  �    9  l  �  �  )  \  �  �  	  G	  }	  �	  �	  .
  `
  �
  �
    >  s  �  �  #  X  �  �     7  l  �  �    S  �  �  �  4  h  �  �  �  ]  ~  �  �  �  �     S  �  �  �  �    ?  �  �  �  /  [  �  �    L  }  �  �  7	  n	  �	  �	  
  Z
  �
  �
  �
  ;  y  �  �    \  �  �    ?  z  �  �  !  Z  �  �  
  D  {  �  �  )  O  i  �  �  �    2  m  �  �  �    N  �  �  �    @  g  �  �    A  o  �  �  	  Q	  �	  �	  �	  *
  f
  �
  �
    B  �  �  �    \  �  �    =  y  �  �  '  \  �  �    D  z  �  �  *  b  �  �  �  �  )  _  �  �  �  *  ^  �  �    +  W  �  �    2  \  �  �  �  -	  ]	  �	  �	  �	  0
  e
  �
  �
  �
  5  l  �  �  	  >  v  �  �    L  �  �  �  )  ]  �  �    =  q  �  �    Q    �  �  �  O  �  �  �    S  �  �  �  (  ^  �  �    @  n  �  �  "	  S	  �	  �	  �	  ,
  b
  �
  �
  �
  6  n  �  �  	  A  z  �  �    I    �  �    S  �  �  �  '  \  �  �  �  0  e  �  z  �  �    V  �  �  �  "  d  �  �    ?  y  �    0  [  �  �  	  K	  y	  �	  �	  *
  d
  �
  �
  �
  ?  |  �  �    W  �  �     6  q  �  �    S  �  �    :  p  �  �    V  �  �  �  1  �  �    �  F  �  �    #  ]  �  �    ;  t  �  �  *  Z  �  �  	  H	  w	  �	  �	  *
  e
  �
  �
  	  H  �  �  �  '  e  �  �    L  �  �  �  6  n  �  �  !  X  �  �    @  x  �  �  #  (  �  �    p  �  �  �    T  �  �  �  !  ]  �  �    3  f  �  �  	  J	  |	  �	  �	  $
  ^
  �
  �
  �
  8  r  �  �    P  �  �  �  -  f  �  �    C  z  �  �  &  \  �  �    =  u  �  �    �    �  �  �    >  �  �  �    @  �  �    9  l  �  �    R  �  �  �  7	  k	  �	  �	  
  R
  �
  �
  �
  4  m  �  �    P  �  �  �  6  o  �  �    S  �  �  �  7  n  �  �    W  �  �  �  T  �  �  �  �  D  �  �    '  [  �  �  "  E  r  �  �  7  c  �  �  	  N	  	  �	  �	  )
  e
  �
  �
    A  ~  �  �    Z  �  �    9  t  �  �  !  V  �  �    =  s  �  �  !  Y  �  �  3  '  �  �    O  Z  �  �    S  }  �  �    R  �  �  �  &  Z  �  �  �  6	  i	  �	  �	  
  J
  
  �
  �
  &  `  �  �     ;  w  �  �    R  �  �  �  1  j  �  �    L  �  �  �  1  g  �  �    ]  �  �  "  q  �  �  �  �  E  {  �  �    ?  �  �  �  &  [  �  �  	  K	  	  �	  

  D
  s
  �
  �
  +  g  �  �    J  �  �  �  +  j  �  �    N  �  �     7  p  �  �    W  �  �  m  ^  q  �  ]  �  �  )  u  �  �  �  7  �  �    5  }  �  �  .  j  �  �  -	  ]	  �	  �	  
  N
  �
  �
  �
  8  m  �  �    W  �  �    >  x  �  �  $  ]  �  �    =  v  �  �    W  �  �  �  n  u  c  q  �  �  �  f  �  �  �  M  �  �  �  8  |  �  �  *  a  �  �  
	  ?	  |	  �	  �	  $
  ]
  �
  �
    G  �  �  �  '  `  �  �    7  h  �  �    J  �  �  �  1  i  �  �    P  �  5  �  �  �    |  �  �  T  �  �  �  '  m  �  �  	  :  v  �  �    D  z  �  �  ,	  a	  �	  �	  
  N
  �
  �
  �
  5  t  �  �     ^  �  �    J  �  �     :  v  �  �  .  i  �  �     ]  �  /  �  �  �  B  v  �  �    a  }  �  �    A  �  �  �  2  g  �  �  1  f  �  �  2	  g	  �	  �	  '
  h
  �
  �
    _  �  �    V  �  �    W  �  �    Q  �  �    F  �  �  �  8  t  �  �  0  �  �  �  4  ~  s  �  �  �  6  �  �  �  ,  }  �    7  y  �    C  {  �  
	  I	  �	  �	  
  K
  �
  �
    G  �  �    D  �  �    ?  �  �    >  {  �  �  :  u  �  �  0  l  �  �  $  /  w  X    �  �  )  �  �  �    r  �  �    ]  �  �    V  �  �  &  Y  �  �  *	  c	  �	  �	  &
  f
  �
  �
  !  c  �  �    ]  �  �    U  �  �    L  �  �    B  �  �  �  8  |  �  �  @  _  .  [  �  �  �  Z  �  �  �  <  �  �  �  !  n  �  �  "  ]  �  �  $  [  �  �  	  Q	  �	  �	  
  K
  �
  �
    ?  {  �  �  -  i  �  �    R  �  �    M  �  �    D  }  �  �  /  e  X  �    >  s  �  �    _  �  �  �  6  }  �  �    `  �  �    H  �  �  �  5  g  �  �  	  J	  �	  �	  
  7
  o
  �
  �
    Q  �  �  �  5  x  �  �    Z  �  �    >  x  �  �    W  �  n  m  �    ;  u  �  �     H  �  �  �    H  �  �  �    R  �  �  �    ]  �  �  �  +  f  �  �  	  9	  q	  �	  �	  
  E
  |
  �
  �
     R  �  �  �  ,  _  �  �    8  k  �  �    C  w  �  d  b  �    :  b  �  �  �    K  �  �  �  �  F  �  �  �    >    �  �  #  L  �  �     1  ]  �  �  	  :	  l	  �	  �	  
  C
  y
  �
  �
    J  �  �  �    R  �  �  �  '  [  �  �  �    Y  `  [  �  �    L  �  �  �    I  �  �  �  �  ;  �  �  �  
  0  y  �  �    A  k  �  �  (  U  z  �  �  (	  \	  �	  �	  �	  *
  d
  �
  �
  �
  (  a  �  �  �  *  ^  �  �    1  `  �  �  �  0  U  �  z  �     M  �  �  �  �  5  p  �  �  �    `  �  �  �    F  �  �    (  :  w  �  �  5  U  k  �  �  -	  a	  �	  �	  �	   
  \
  �
  �
  �
    P  �  �  �  �  <    �  �  
  �  �    O  �  |  h  �    p  �  �  �    d  �  �  �    W  �  �  �    C  �  �  �    A  z  �  �    B  o  �  �  	  H	  p	  �	  �	  
  I
  r
  �
  �
    F  s  �  �    =  r  �  �    ,  b  �    z  �  q  �     _    �  �    T  �  �  �  �  ;  s  �  �  �  !  Z  �  �  �    F  �  �  �    7  o  �  �  �  )	  `	  �	  �	  
  )
  W
  �
  �
    ,  U  �  �  �  ,  R  }  �  ,  .  �  �  s  w  q  �  �  F  X  �  �  �    C  [  ~  �  �  '  K  k  �  �    @  d  �  �  �  6  e  �  �  �  $  a  �  �  �  	  P	  �	  �	  �	  
  B
  �
  �
  �
    9  w  �  �    >  n  �  r  �        j  �  �    /  9  I  n  �  �  �    K  �  �  �    =  v  �      =  r  �  �  /  <  l  �  �  +  X  i  �  �   	  ^	  �	  �	  �	  
  Y
  �
  �
  �
    O  �  �  �    I  �  �    h  A  v  |  �  �  �  �  �  �  >  y  �  �  �    ^  �  �  �    I  �  �  �    D  �  �  
  /  S  �  �    @  c  �  �  	  J	  t	  �	  �	  
  I
  �
  �
  �
    E  �  �  �    C    4  P  �  b  a  �  �  �  �  �  �  �  &  O  �  �  �  �  V  �  �  �  �  C  �  �  �    <  �  �    '  G  �  �    B  `  �  �  	  R	  y	  �	  �	  
  Y
  �
  �
  �
    Y  �  �  �    V  Y  d  X  f  �  �      '  4  F  j  �  �  �  �  �    U  �  �  �  �  -  |  �  �  �  %  p  �  �    4  h  �  �  ,  N  r  �  �  9	  f	  �	  �	  �	  >
  w
  �
  �
  �
  =  |  �  �    =    c  c  �  �    ,  \  ~  �  �  �  �    :  b  �  �  �  �    D  o  �  �  �  �  '  [  �  �    *  R  �  �    9  ]  �  �  	  E	  o	  �	  �	  
  M
  �
  �
  �
  
  K  �  �  �    N  �  �  X  �  �  0  V  {  �  �  �  !  H    �  �  �    G  z  �  �     #  T  �  �  �    9  b    �  �  
  B  w  �  �  	  9	  o	  �	  �	  �	  /
  m
  �
  �
  �
  .  i  �  �    5  l  �  �    B  y  �    U  �  �  �    V  �  �  �    <  s  �  �    B  r  �  �    9  c  �  �    4  R  �  �  �  #	  W	  �	  �	  �	  
  L
  �
  �
  �
    O  �  �  �  !  Y  �  �  �  "  S  �  �  �  �  �    S    �  �  *  h  �  �  �  3  w  �  �  
  A  z  �  �  "  c  �  �    :  v  �  �  	  T	  y	  �	  �	  
  U
  �
  �
  �
  /  Z  �  �    ;  s  �  �    M  �  �  �  ,  O  �  �  �  �  �  *  a  �  �    \  �  �  �  -  �  �  �    [  �  �  	  A  z  �  �  3  z  �  �  -	  d	  �	  �	  
  L
  �
  �
  �
  #  j  �  �    J    �  �  ,  f  �  �    G  }  �  �  &  ^  |  |  |  K  �  �  �  �    g  �  �    g  �  �    @  �  �    :  {  �  �  6  m  �  �  )	  e	  �	  �	  
  `
  �
  �
    N  �  �    9  r  �  �  #  [  �  �    G  �  �  �  0  o  �  �    !  !  k  �  �  �  �    o  �  �  
  ^  �  �    K  �  �    B  �  �    D  w  �   	  >	  s	  �	  �	  ,
  k
  �
  �
    \  �  �    M  �  �    @  {  �  �  0  i  �  �    X  �  �    G  �  �  r  �  �  ,  {  W  �  �  �  �  D  �  �  �  -  s  �  �  %  ]  �  �  %  V  �  �  	  Q	  �	  �	  
  C
  }
  �
  �
  *  k  �  �    U  �  �    E  �  �  �  :  s  �  �  *  c  �  �    P  �  �  �  �  B  �  �  �  �  3  �  �  �  �  )  e  �  �    2  g  �  �    E  x  �  �  *	  ^	  �	  �	  
  D
  z
  �
  �
  #  `  �  �    B    �  �  (  c  �  �    L  �  �  �  9  r  �  �  !  �  �  �  ?  �  �  �  �  7  �  �  �    H  �  �  
  3  `  �  �    I  u  �  �  &	  \	  �	  �	  �	  3
  n
  �
  �
    C  �  �  �    W  �  �  �  .  e  �  �    @  v  �  �    S  �  �  �  �  �  �  $  s  �  �    b  �  �    ?  v  �  �  '  X  �  �    @  s  �  �  #	  ]	  �	  �	  
  @
  z
  �
  �
  $  _  �  �  
  D    �  �  +  e  �  �    I  �  �  �  -  g  �  �    K  �    !  k  6  v  �    2  a  �  �    7  l  �  �  %  U  �  �    M  �  �  	  @	  t	  �	  �	  *
  f
  �
  �
    J  �  �  �  5  q  �  �  $  ^  �  �    I  �  �  �  3  k  �  �    T  �  �  �  B  �  �  �  �    G  �  �  	  =  u  �  �    I  �  �  �  ,  ]  �  �  	  F	  z	  �	  �	  -
  f
  �
  �
    B  �  �  �  .  f  �  �    A  y  �  �  #  [  �  �  	  A  w  �  �  !  Z  �  �    J  �  �     5  �  �  �    ;    �  �  /  f  �  �    I  �  �  �  -	  b	  �	  �	  
  H
  ~
  �
  �
  +  d  �  �    G  �  �  �  -  f  �  �    J  �  �  �  /  f  �  �    O  �  �  �  )  �  �  �  �  6  ~  �    $  R  �  �    @  k  �  �  +  \  �  �  	  A	  w	  �	  �	  
  X
  �
  �
  �
  5  q  �  �    O  �  �  �  1  j  �  �    M  �  �  �  3  j  �  �    O  �  �  �  "  r  �  �  7  A  k  �    A  `  �  �  �  :  n  �  �  �  6  r  �  �  	  ;	  x	  �	  �	  
  L
  �
  �
  �
  ,  a  �  �    D  y  �  �  &  \  �  �    =  u  �  �    V  �  �  �  6  p  @    	  P  �    0  @  s  w  �    A  k  �  �    I  {  �  �  *  c  �  �  	  M	  �	  �	  �	  7
  v
  �
  �
  &  a  �  �    K  �  �  �  3  o  �  �     X  �  �    E  }  �  �  0  i  �  1  �    g  	  P  �  �    M  �  �  �  >  �  �    8  {  �  �  ?  v  �  �  4	  q	  �	  �	   
  \
  �
  �
    C  �  �  �  '  e  �  �    O  �  �    <  u  �  �  *  a  �  �    L  �  �  �  
  ,  �    M  �  �     U  �  �    M  �  �    K  �  �    A  w  �  �   	  U	  �	  �	  �	  @
  x
  �
  �
    a  �  �  
  G  �  �  �  1  m  �  �    R  �  �  �  8  p  �  �    V  �  �  �  �  �  )  E  �  �  �  B  �  �  �  9  m  �  �    O  �  �    K    �  �  5	  l	  �	  �	  
  V
  �
  �
  �
  :  }  �  �  &  d  �  �    Q  �  �  
  C  ~  �  �  7  q  �  �  (  e  �  �  V  s  �  �  '  [  �  �    X  �  �    @  �  �     9  h  �  �  3  k  �  �  1	  n	  �	  �	  (
  e
  �
  �
    W  �  �    F  �  �  �  ;  z  �  �  3  o  �  �  ,  h  �  �  #  a  �  �  �    V  �  �    4  g  �  �    X  �  �    E  }  �  �  ?  {  �  �  ?  }  �  �  ;	  z	  �	  �	  :
  x
  �
  �
  6  s  �  �  0  m  �  �  (  g  �  �  "  `  �  �    [  �  �    W  �  �  �  �  9  ~  �  �  �  -  Q  �  �    A  �  �  	  D  }  �    B  {  �  �  >  z  �  �  <	  z	  �	  �	  9
  z
  �
  �
  7  w  �  �  4  s  �  �  .  m  �  �  %  b  �  �    X  �  �    W  �  �    �  '  2  �  �  �    P  �  �  
  C  �  �  	  B  �  �    >  ~  �  �  8  u  �  �  ,	  l	  �	  �	  %
  `
  �
  �
    T  �  �    @  y  �  �  #  c  �  �    S  �  �  �  8  g  �  �  X  X  �  �    *  v  �  �    O  �  �  	  C    �  �  3  m  �  �     X  �  �    ?  ~  �  �  "	  i	  �	  �	  
  G
  �
  �
  �
    N  �  �  �  (  [  �  �  �  (  \  �  �  �  2  g  �  �  n  Y  Z  �  �  �     x  �  �    ;  z  �  �    K  �  �  �  )  \  �  �    8  k  �  �    F  z  �  �  	  Q	  �	  �	  �	  
  Z
  �
  �
  �
  *  c  �  �    7  m  �  �    D  x  �  �    �  �  W  X  �  �  �    N  �  �  �    [  �  �  �    [  �  �  �  &  a  �  �    7  h  �  �    E  q  �  �  	  T	  �	  �	  �	  "
  [
  �
  �
  �
  (  `  �  �  �  .  e  �  �  �  3  i  �  �  �  �    X  a  �  �  7  b  �  �  �  !  m  �  �  �    _  �  �  �  !  V  �  �  �  $  Z  �  �     *  Y  �  �  �  (	  X	  �	  �	  �	  ,
  ^
  �
  �
  �
  *  ^  �  �  �  (  Z  �  �  �  $  �  �  �    ]  j  �  �  �  7  y  �  �  �    `  �  �  �  �  3  |  �  �  �    V  �  �  �    F  �  �  �    E  q  �  �  	  =	  n	  �	  �	  

  7
  e
  �
  �
  �
  1  _  �  �  �  (  Y  �  ,  L  �  �  +  g  a  v  �     >  T  �  �  �  �  (  [  �  �  �    ;  l  �  �    :  _  �  �    =  _  �  �  �  <  k  �  �  �  /	  m	  �	  �	  �	  !
  c
  �
  �
  �
    U  �  �  �    O  ,  ,  ,  �    P  \  q  �  �  �  �    F  �  �  �  �  -  u  �  �  �    c  �  �      E  �  �    /  9  n  �    C  ]  p  �  �  =	  t	  �	  �	  �	  .
  q
  �
  �
  �
    f  �  �  �    ,  .  �  �        �  $  v  �  �  �  �  T  �  �  �  �  8  �  �  �  �  .  |  �  �  
  4  q  �  �  %  >  i  �  �  1  T  o  �  �  /	  f	  �	  �	  �	  &
  i
  �
  �
  �
    c  �  �  �    �  r  �  V  @  >  z  j  �    �  �  �  �    j  �  �  �    _  �  �  �    T  �  �  �    R  �  �    3  Z  �  �  #  K  k  �  �  %	  \	  �	  �	  �	  #
  e
  �
  �
  �
    d  �  �  �  !  �  �    -  �  �  �  �  �     k  h  n  �  )  m  �  �  �    f  �  �  �  
  Y  �  �  �    R  �  �    -  W  �  �  #  H  j  �  �  +	  ^	  �	  �	  �	  +
  j
  �
  �
  �
  *  n  �  �  �  -    4  K  )       8  E  X  p  �  �  �    I  �  �  �  �  >  �  �  �  �  .  �  �  �  �  '  u  �  �    7  q  �    6  S  z  �  		  G	  n	  �	  �	  
  M
  �
  �
  �
    N  �  �  �    O  >  Y  X  f  p  y  |  �  �  �    L  v  �  �  �    :  l  �  �  �    G  �  �  �  	  9  �  �  �     C  v  �    1  T  ~  �  	  @	  j	  �	  �	  
  H
  }
  �
  �
  
  I  �  �  �    K  �  X  c  p  v  �  �  �  .  V  q  �  �  �    =  }  �  �  �  8  i  �  �  �    K  �  �  �    D  s  �  �    L  |  �  �  		  I	  �	  �	  �	  
  R
  �
  �
  �
    P  �  �  �  '  Y  �  �  �  X  �  �  �  �  #  c  }  �  �  �  )  a  �  �  �  "  Z  �  �    2  d  �  �    A  o  �  �    6  k  �  �  	  <	  u	  �	  �	  
  I
  �
  �
  �
    S  �  �  �  0  h  �  �    7  i  �  �  y  �    R  Q  s  �  �  �  /  t  �  �  �  9  x  �  �    C  �  �  �  )  `  �  �    ?  v  �  �  	  O	  �	  �	  �	  7
  o
  �
  �
    L  �  �  �  /  e  �  �    D  {  �  �    S  �  �  �    R  y  �  �  �  �  8  �  �  �  #  `  �  �    I  �  �  �  3  n  �  �    Q  �  �  	  ;	  r	  �	  �	  &
  [
  �
  �
    E  �  �  �  5  p  �  �    T  �  �    ?  {  �  �  )  ]  ]  �  *  Y  �  �  �    :  ~  �  �    d  �  �    Q  �  �    H  �  �    M  �  �  	  A	  x	  �	  �	  4
  m
  �
  �
    b  �  �    P  �  �  �  ;  z  �  �  .  j  �  �    T  �  �      J  y  n  �  �    c  �  �  �  	  ?  �  �  �  1  z  �  �  6  u  �  �  8  r  �  �  9	  x	  �	  �	  7
  t
  �
  �
  *  j  �  �     _  �  �    S  �  �    J  �  �    ?  }  �  �  1  n  q  e  �  �  �  �    l  �  �  �  5  }  �  �  	  E  �  �    4  t  �  �  7  n  �  �  5	  n	  �	  �	  .
  o
  �
  �
  '  i  �  �    _  �  �    U  �  �    L  �  �    C  �  �  �  :  v  �  h  �  �  (  s  U  �  �  �  �  A  �  �  �    Z  �  �    5  o  �  �  )  W  �  �  	  N	  �	  �	  �	  =
  y
  �
  �
  &  h  �  �    W  �  �    K  �  �    A  ~  �  �  5  m  �  �  &  a    �  �  >  �  �  �  �  /  �  �  �  �  !  b  �  �  �  '  ^  �  �    5  f  �  �  	  I	  y	  �	  �	  $
  ]
  �
  �
  �
  9  u  �  �    R  �  �  �  6  q  �  �  !  Y  �  �    F    �  �  �  �  �  =    �  �  �  4  �  �  �    D  �  �     )  Z  �  �    ?  m  �  �  	  R	  �	  �	  �	  +
  c
  �
  �
  �
  :  t  �  �    L    �  �     W  �  �  �  /  e  �  �  	  ?  u  �  �  �  �  �  "  m  �  �    _  �  �  �  8  q  �  �    O  �  �  �  5  j  �  �  	  S	  �	  �	  �	  8
  q
  �
  �
    X  �  �    <  w  �  �  #  ]  �  �    A  z  �  �  %  _  �  �    C  }  
    c  &  j  �    -  Y  �  �    0  g  �  �    M  �  �    C  {  �  �  7	  k	  �	  �	  #
  ]
  �
  �
  
  C  }  �  �  -  j  �  �    V  �  �    A  z  �  �  *  c  �  �    K  �  �  �  @  y  �  �  �  �  D  �  �  �  6  p  �  �    A  }  �  �  $  T  �  �  	  >	  q	  �	  �	  %
  ]
  �
  �
     9  z  �  �  %  ^  �  �    9  q  �  �    R  �  �    9  o  �  �    Q  �  -  P  �  6  `  �  �  9    U  �  �  1  ]  �  �  #  T  �  �    S  �  �  
	  O	  �	  �	  �	  ?
  �
  �
  �
  ,  s  �  �     _  �  �    T  �  �    N  �  �    A  {  �  �  8  r  �  �  $  +  n  �    q  �  �  �  5  z  �  �    F  �  �  �  6  l  �  �    X  �  �  	  G	  }	  �	  �	  4
  m
  �
  �
    V  �  �  �  5  y  �  �  "  \  �  �    H  �  �  �  5  p  �  �  $  ^  �  d  �  �  �  2  u  �  �  �  :  |  �  �  �  9  |  �  �  	  :  w  �  �    C  z  �  �  (	  X	  �	  �	  
  ;
  o
  �
  �
    O  �  �  �  *  e  �  �  	  B  ~  �  �  &  ^  �  �    D  |  �  t  �  O  �  %  ,  f  {  �  �  �  M  m  �  �  �  ;  x  �  �    R  �  �    C  y  �  	  ;	  p	  �	  �	  .
  j
  �
  �
    Y  �  �  
  I  �  �  �  ;  z  �  �  2  n  �  �  *  f  �  �     i  )  F  �  O  �      O  �  �  �  /  �  �  �  %  q  �  �  /  j  �     6  k  �  �  :	  p	  �	  �	  2
  t
  �
  �
  *  p  �  �  $  f  �  �  %  a  �  �  #  `  �  �  "  _  �  �    _  �  �  5  i  *  @  �  �  �  T  �  �  �  A  �  �  �  @  �  �    C  �  �    K  �  �  	  S	  �	  �	  
  U
  �
  �
    Q  �  �    N  �  �    N  �  �    O  �  �    P  �  �    R  �  �  4  �  �  �  [  z  �  �  A  �  �  �  0  �  �  �  '  s  �  �  0  o  �  �  8  q  �  �  9	  t	  �	  �	  7
  v
  �
  �
  2  u  �  �  /  q  �  �  .  n  �  �  .  m  �  �  .  l  �  �  -  l  �  $  �  z  �  5  i  �  �    d  �  �  �  B  �  �  �  /  v  �  �  +  f  �  �  *  f  �  �  ,	  g	  �	  �	  *
  h
  �
  �
  &  h  �  �  #  f  �  �  #  d  �  �  #  c  �  �  $  c  �  �  (  g    X  Z  �  �  L  k  �  �    ^  �  �  �  >  �  �  �  .  z  �  �  1  u  �  �  5  r  �  �  :	  v	  �	  �	  ;
  z
  �
  �
  ;  |  �  �  :  |  �  �  9  {  �  �  8  y  �  �  7  v  �  �  4  �  ?  ^  �  �  �  9  r  �  �    S  �  �  �  A  �  �  �  8  �  �  �  5  x  �     ;  y  �  �  <	  y	  �	  �	  :
  x
  �
  �
  5  s  �  �  .  l  �  �  %  b  �  �    X  �  �    R  �  �    3  !  �  Z  �  �  -  a  �  �    W  �  �    K  �  �  �  <  �  �  �  8  w  �  �  +  i  �  �  #	  `	  �	  �	  
  R
  �
  �
    >  w  �  �  &  ]  �  �  !  X  �  �    O  �  �    ;  ,  �      F  [  �  �  &  a  �  �    L  �  �  �  :  t  �  �  "  X  �  �    <  s  �  �    U  �  �  	  B	  |	  �	  �	  #
  \
  �
  �
    K  �  �  �  )  f  �  �    E  z  �  �  #  W  �  ,  �  �    ;  f  �  �    L  y  �  �    [  �  �  �  (  b  �  �  �  2  k  �  �  �  7  t  �  �    =  {  �  �  	  D	  �	  �	  �	  
  N
  �
  �
  �
  +  Z  �  �    6  f  �  �  	  @  �  ,  ,  `  �  	  C  J  d  �    &  F  n  �  �    >  r  �  �  	  +  s  �  �    8  k  �  �  &  L  q  �  �  ,  `  �  �  �  0	  k	  �	  �	  �	  3
  q
  �
  �
    9  s  �  �    C  x  �  ,  ,  ,  2  �  �  �  �  7  w  �  |  �  /  u  �  �  �  %  d  �  �  �    Y  �  �      P  �  �    <  [  �  �    H  r  �  �  	  P	  �	  �	  �	  
  J
  �
  �
  �
    ?  �  �  �    E  �   �   �   4  �  B  8  �  �  9  �  �  o  �    Y  �  �  �  �  ;  �  �  �  �  &  o  �  �      Z  �  �  +  3  C  �  �  #  X  c  {  �  	  V	  �	  �	  �	   
  H
  �
  �
  �
  �
  9    �  �  �  �   �   �   "  �  H  ,  �  �  U  �  }  �  �  O  �  �  �  �  B  �  �  �  �  7  �  �  �    9  �  �    *  G    �    D  _  �  �  	  O	  y	  �	  �	  
  N
  �
  �
  �
  �
  ;  �  �  �                �   �   �  �  l  �  �  q  t  x  �  �  [  �  �  �  �  S  �  �  �  �  H  �  �  �  	  >  �  �    *  F  �  �    D  `  �  �  	  P	  y	  �	  �	  

  P
  �
  �
  �
    J  �  �  �                �   �   �  L  K  �  �  J  s  {  �  �  I  �  �  �  �  @  �  �  �  �  9  �  �  �    :  �  �  	  '  H  �  �    A  _  �  �  	  S	  y	  �	  �	  
  Z
  �
  �
  �
    W  �  �  �    �  �   �   �      y  ,  6  �  �  H  �  d  �  �  E  �  �  �  �  ?  �  �  �  �  5  �  �  �    7  �  �    #  E  �  �    >  ]  �  �  	  R	  w	  �	  �	  
  [
  �
  �
  �
    ]  �  �  �    �   �   �   6  ?  ,  �  �  �     f  \  ]  �  "  _  �  �  �  	  \  �  �  �  �  P  �  �  �    F  �  �    #  L  �  �    ?  _  �  �   	  T	  x	  �	  �	  !
  a
  �
  �
  �
  "  f  �  �  �  (  N  V  |  0  R  �  �  "  X  f  �  �  �  0  _  �  �  �    Z  �  �  �    P  �  �  �    F  �  �    '  M  �  �    C  b  �  �  &	  Y	  |	  �	  �	  (
  h
  �
  �
  �
  +  p  �  �  �  1  r  �  ,  ,  g  �  �  8  h  y  �  �  H  t  �  �  �  ?  {  �  �  �  2  i  �  �    3  d  �  �    H  y  �  �    J  |  �  �  	  Y	  �	  �	  �	  ,
  h
  �
  �
    5  m  �  �    .  _  �  �  F  W  �  �    N  x  w  �  $  W  �  �  �  -  x  �  �    Q  �  �  �  )  _  �  �    7  u  �  �    T  �  �  �  )	  g	  �	  �	  
  K
  �
  �
  �
  .  e  �  �     6  h  �  �  �  0  _  �  ,  �  �  5  s  q  �  �    [  �  �  �  I  �  �  �  &  j  �  �    Q  �  �    E  �  �  �  0  h  �  �  	  L	  �	  �	  
  <
  u
  �
  �
  '  _  �  �    G  �  �  �  +  b  �  �    K    ~  �    i  e  �    G  �  �  �    X  �  �  �  3  w  �  �    ]  �  �    O  �  �    D  ~  �  �  6	  t	  �	  �	  ,
  h
  �
  �
     \  �  �    L  �  �  �  :  w  �  �  '  c  �  �    )     ^  ~  �  �  <  �  �  �    q  �  �  �  M  �  �  �  -  y  �  �  $  \  �  �  &  W  �  �  	  V	  �	  �	  
  L
  �
  �
  �
  >  }  �  �  /  p  �  �  #  b  �  �    U  �  �    J  �  b    �  q  �  +  h  �  �    `  �  �    T  �  �    B  �  �    <  �  �    D  �  �  	  E	  �	  �	  
  B
  �
  �
    A  �  �  �  8  x  �  �  :  x  �  �  6  r  �  �  .  j  �  �  3  �  �  �  q  �  ,  q  �  �  !  z  �  �    m  �  �    h  �  �  ,  i  �  �  6  k  �  �  <	  q	  �	  �	  8
  t
  �
  �
  4  w  �  �  4  u  �  �  1  p  �  �  4  s  �  �  4  s  �  �  1  p  k  �  ,  r    @  ~  �  �  %  q  �  �    d  �  �    T  �  �  &  X  �  �  .  b  �  �  ,	  h	  �	  �	  *
  j
  �
  �
  !  f  �  �    `  �  �    ]  �  �    Z  �  �    X  �  �    V  e  �  9  e  �  �  �  %  6  ?  q  �  �    Q  �  �    .  x  �  �  -  c  �  �  -  _  �  �  &	  a	  �	  �	  
  U
  �
  �
    K  �  �    C  �  �  �  <  |  �  �  6  v  �  �  )  f  �  �    ?  �  �  �  �  �  [  �  �  �    O  �  �  �    A  {  �  �  
  ?  w  �  �    P  �  �  �  4	  h	  �	  �	  
  O
  �
  �
  �
  2  n  �  �    T  �  �    ?  z  �  �  .  i  �  �    V  �  5  m  �  �    F  �  �     7  j  �  �    O  �  �  �  '  \  �  �    9  l  �  �  	  I	  	  �	  �	  #
  [
  �
  �
     7  n  �  �    <  s  �  �    E  {  �  �  !  S  �  �  �  .  b  �  s  �  �  ,  }  �  �  �  ,  �  �    #  X  �  �    R  �  �    <  |  �  �  2	  n	  �	  �	  
  Y
  �
  �
  �
  6  s  �  �  $  ^  �  �    E  �  �  �  +  d  �  �    <  r  �  �  )  _  �    �  �  
  r  �  �  
  S  �  �    R  �  �     J  �  �    S  �  �  	  G	  	  �	  �	  :
  x
  �
  �
  *  e  �  �    Z  �  �    K  �  �  �  4  n  �  �  *  c  �  �    J  �  �  �  �  $  �    $  g  �  �  4  �  �    "  U  �  �  ,  a  �  �  1  c  �  �  &	  f	  �	  �	  
  [
  �
  �
    L  �  �    B  �  �  �  8  v  �  �  /  j  �  �     \  �  �    <  t  �  �    2  ]  �  8  h  �  �  8    P  �  �  /  X  �  �    Q  �  �    L  �  �  �  E	  }	  �	  �	  4
  x
  �
  �
  #  h  �  �    V  �  �    M  �  �    F  �  �  �  =  x  �  �  /  l  �  �    /    �    �  �  �  �  5  �  �  �    F  �  �  �  ;  l  �  �  !  [  �  �  	  F	  	  �	  �	  0
  m
  �
  �
    Q  �  �  �  6  t  �  �  "  [  �  �    I  �  �  �  8  q  �  �  #  _  �  �  �  �  �  0  �  �  �  �  7  �  �  �    :  �  �  �    ?  |  �  �    K  �  �  �  1	  a	  �	  �	  
  C
  x
  �
  �
    W  �  �  �  0  l  �  �    J  �  �  �  /  f  �  �    M  �  �  �  �  ]  �    5  j  �  �  �    L  t  �  �    =  z  �  �  +  W  �  �    P    �  	  G	  {	  �	  �	  5
  u
  �
  �
    `  �  �    O  �  �    C  �  �     ;  v  �  �  2  o  �  �  )  x  *  [  �  \  �    "  O  �  �  �  .  �  �    %  s  �    9  k  �    D  s  �  �  F	  |	  �	  �	  :
  
  �
  �
  0  y  �  �  +  m  �  �  -  i  �  �  -  i  �  �  +  i  �  �  '  g  �  �  5  �  *  N  �  �  �  V  �  �  �  B  �  �    @  �  �    I  �  �     V  �  �  	  ^	  �	  �	  
  `
  �
  �
    Z  �  �    V  �  �    V  �  �    W  �  �    X  �  �    [  �  �  D  �  �  �  c  �  �  �  E  �  �  �  0  �  �  �  +  w  �    9  s  �    C  x  �   	  D	  ~	  �	  �	  @
  �
  �
  �
  :  ~  �  �  7  z  �  �  6  w  �  �  7  u  �  �  7  u  �  �  6  u  �  1  �  u  �  7  �  �  �    o  �  �  �  D  �  �    3  {  �    4  l  �  �  5  n  �  �  7	  q	  �	  �	  2
  s
  �
  �
  -  q  �  �  +  m  �  �  +  k  �  �  ,  j  �  �  ,  j  �  �  /  n    �  \  �  �  _  ~  �  �    c  �  �  �  @  �  �  �  3    �    ;  z  �    A  {  �  	  E	  �	  �	   
  D
  �
  �
  �
  B  �  �     @  �  �  �  =  ~  �  �  <  {  �  �  9  v  �  �  /  �  `  r  �  �  �  =  �  �  �    [  �  �  �  E  �  �    =  �  �    >  ~  �    E  �  �  	  F	  �	  �	   
  A
  ~
  �
  �
  6  t  �  �  %  d  �  �    O  �  �  �  :  t  �  �  &  Z  Z    2  .  �  g  �  �  5  y  �  �    `  �  �    O  �  �    A  �  �    >  |  �  �  /  i  �  �  	  X	  �	  �	  �	  5
  m
  �
  �
    A  w  �  �    T  �  �  �  1  h  �  �    4  h  �  ,  �      h  k  �  �  +  p  �  �    R  �  �  �  >  |  �  �  '  ^  �  �    #  [  �  �  �    I  �  �  �  	  K	  |	  �	  �	  
  J
  �
  �
  �
  (  T  {  �  �  %  V  �  �  �  -  `  �  x  ,  �  �    O  i  �  �    X  �  �  �  "  a  �  �  �  ,  ]  �  �  �  '  I  c  �  �    I  k  �  �    N  {  �  �  	  F	  	  �	  �	  
  I
  �
  �
  �
    O  �  �  �    O  �  �  �  �  ,  ,  `  �  	  `  g  j  �    +  S  v  �  �    ?  w  �  �  �  %  h  �  �    /  W  �  �    ?  b  �  �    <  k  �  �  �  2	  l	  �	  �	  �	  ,
  l
  �
  �
    ,  c  �  �    6  Z  G  v  Z  2  �  �  �  �  7  w  �  z  �  /  v  �  �  �    L  �  �  �  �  6  �  �       '  n  �    /  A  d  �  �  :  `  y  �  �  )	  g	  �	  �	  �	  
  _
  �
  �
  �
     F  �  �  �    �   �   �   4  �  B  8  �  �  9  �  x  m  �    Y  �  �  �  �  :  �  �  �  �    k  �  �  �    N  �  �  "  *  ;  �  �    O  Z  r  �  
	  N	  ~	  �	  �	  �	  A
  �
  �
  �
  �
  /  x  �  �  �  �   �   �   "  �  E  ,  �  �  R  �  |  �  �  E  �  �  �  �  6  �  �  �  �  (  �  �  �    +  t  �  �    =  s  �    7  V  |  �  	  D	  o	  �	  �	   
  G
  
  �
  �
  �
  :  �  �  �  �              �   �   �  �  l  �  �  L  c  b  �  �  G  �  �  �  �  >  �  �  �  �  6  �  �  �    8  �  �    $  F  �  �    @  _  �  �  	  R	  x	  �	  �	  
  W
  �
  �
  �
    T  �  �  �                �   �   j  3  ,  �  �  D  y  e  �  �  C  �  �  �  �  >  �  �  �  �  5  �  �  �     4  �  �      A  �  �    ;  Y  �  �  	  O	  s	  �	  �	  
  Z
  �
  �
  �
    ^  �  �  �    g  �   �   �      s  ,  6  �  �  i  s  \  �    \  �  �  �     Z  �  �  �    W  �  �  �    U  �  �    +  \  �  �  )  I  m  �  �  7	  c	  �	  �	  �	  @
  x
  �
  �
     F  �  �  �    L  �   �   �   6  >  ,  �  �    G  [  t  �    @  q  �  �  �  1  u  �  �  �  %  q  �  �  �  '  i  �  �    8  j  �  �  +  O  v  �  �  8	  e	  �	  �	  �	  >
  v
  �
  �
  �
  A  �  �  �    F  8  V  ,  0  R  �  �  "  Z  h  �  �  D  r  �  �    F  |  �  �    I  �  �  �  0  ^  �  �    F  s  �  �  $  ^  �  �  �  7	  v	  �	  �	  
  =
  x
  �
  �
    B  t  �  �    L  {  �  �  �  ,  ,  `  �  �  8  [  x  �  $  T  {  �  �  2  q  �  �    E  �  �  �  )  i  �  �    J  �  �  �  2  s  �  �  	  W	  �	  �	  
  >
  z
  �
  �
  %  X  �  �  �  $  Q  x  �  �    G  }  D  P  �  �    ?  U  v  �  "  V    �  �  M  �  �  �  "  o  �  �  	  L  �  �    ;  ~  �  �  3  k  �  �  )	  _	  �	  �	  
  T
  �
  �
    F  ~  �  �  1  o  �  �    M  �  �  �    D  ,  �  �  4  X  g  �  �    R  |  �  �  F  �  �  �  *  y  �  �    a  �  �    S  �  �    K  �  �  	  E	  ~	  �	  
  B
  |
  �
  �
  9  v  �  �  ,  k  �  �    ]  �  �    N  �  �    ~  �    ]  c  �    F  w  �  �    S  �  �  �  /  s  �  �    [  �  �    K  �  �    D  �  �  	  @	  {	  �	  �	  =
  x
  �
  �
  6  u  �  �  -  n  �  �  %  e  �  �    \  �  �    S    �  Q  \  |  �  7  r  �  �    k  �  �  �  H  �  �  �  '  s  �  �    V  �  �    O  �  �  	  N	  �	  �	  
  G
  �
  �
  �
  ;  z  �  �  .  p  �  �  #  d  �  �    Y  �  �    Q  �  <    �  n  �  (  a  �  �    ^  �  �  �  Q  �  �  �  <  �  �    4  ~  �    ;  {  �   	  =	  }	  �	  �	  <
  z
  �
  �
  ;  |  �  �  4  t  �  �  7  u  �  �  5  p  �  �  /  k  �  �  5  ~  �  �  n  �  ,  i  �  �    s  �  �    j  �  �    e  �  �  #  c  �  �  +  c  �  �  2	  h	  �	  �	  0
  l
  �
  �
  -  p  �  �  -  o  �  �  *  k  �  �  /  n  �  �  1  p  �  �  /  n  j  �  ,  i  �  4  t  �  �  "  n  �  �     `  �  �  
  Q  �  �    Q  �  �  $  Y  �  �  $	  ^	  �	  �	  #
  a
  �
  �
    ^  �  �    Y  �  �    R  �  �    >  y  �  �  8  t  �  �  '  d  �  +  ]  �  �  �     0  4  g  �  �    L  �  �  �  (  s  �  �  #  ]  �  �  "  V  �  �  	  W	  �	  �	  
  N
  �
  �
    D  �  �  �  ;  {  �  �  4  t  �  �  .  k  �  �    Z  �  �    "  h  �  �  �  �  I  �  �  �    F    �  �  �  8  r  �  �    6  o  �  �    F  ~  �  �  +	  _	  �	  �	  
  G
  }
  �
  �
  *  f  �  �    L  �  �  �  7  s  �  �  &  a  �  �    M  �  +  f  �  �    7  �  �  �  /  ^  �  �    H  }  �  �    U  �  �  �  0  d  �  �  	  @	  v	  �	  �	  
  Q
  �
  �
  �
  .  e  �  �  �  3  j  �  �    <  r  �  �    J  }  �  �  %  Y  �  O  �  �  #  g  �  �  �  %  z  �  �    Q  �  �    J  �  �    3  t  �  �  (	  e	  �	  �	  

  O
  �
  �
  �
  -  j  �  �    U  �  �  �  <  {  �  �  "  [  �  �  �  3  i  �  �     V  �  #  �  �    o  �  �    I  �  �    K  �  �    D  {  �    K  ~  �  �  =	  w	  �	  �	  0
  n
  �
  �
  !  [  �  �    P  �  �    A  |  �  �  +  d  �  �  !  Y  �  �    E  �  �  �  �    �       V  �  �  .  x  �  �    O  �  �  %  [  �  �  '  \  �  �  	  ]	  �	  �	  

  Q
  �
  �
    B  �  �  �  :  y  �  �  0  m  �  �  &  a  �  �    S  �  �    K  �  �    ?  �  S  s  �  �  �  P  r  �  �    V  �  �  �  .  f  �  �    N  �  �  		  A	  r	  �	  �	  .
  j
  �
  �
    Z  �  �    E  �  �  �  4  o  �  �    N  �  �  �  4  k  �  �    S  �  �  �  �  )  U  b  �  �  
  T  �  �  �  5  |  �  �    [  �  �    >  x  �  �  /	  `	  �	  �	  
  P
  �
  �
  �
  2  n  �  �    P  �  �  �  2  p  �  �    T  �  �    >  u  �  �  '  _  �  �  �  �    {  �  �  �  !  |  �  �    >  �  �  �  '  T  �  �    ;  h  �  �  !	  R	  �	  �	  �	  5
  l
  �
  �
    K  �  �  �  &  d  �  �  
  C  �  �  �  *  b  �  �    L  �  �  �  6  o  �  �    m  �  �  �    o  �  �  �    c  �  �     2  x  �  �  (  Y  �  �  "	  T	  �	  �	  
  P
  �
  �
  �
  B  �  �  �  )  n  �  �    [  �  �    R  �  �    I  �  �     ?  |  �  �  �  �  �  U  S  q  �  �    o  �  �    S  �  �    @  �  �    K  �  �  	  S	  �	  �	  
  T
  �
  �
    M  �  �    D  �  �    =    �     ;  y  �  �  8  u  �  �  3  r  �  �  ,  l  �  �  �  �  ?  q  �  �    t  �  �    `  �  �    ]  �  �  ,  b  �  �  0	  i	  �	  �	  .
  m
  �
  �
  *  k  �  �  #  f  �  �     b  �  �    _  �  �    \  �  �    T  �  �    R  j  *  t  �  �  &  d  �  �  �  Y  �  �    N  �  �    G  �  �    O  �  �  	  O	  �	  �	  
  I
  �
  �
    G  �  �     >  |  �  �  ;  y  �  �  5  p  �  �  (  g  �  �  #  `  �  �      '  X  �  �  �  J  �  �  �  +  w  �  �    Z  �  �    K  �  �  
  @  y  �  �  9	  t	  �	  �	  +
  k
  �
  �
    ^  �  �    O  �  �    @  |  �  �  .  i  �  �    V  �  �    M  y  y  !  ;  s  �  �    S  �  �  �  )  t  �  �    ?  �  �  �  ,  e  �  �     [  �  �  	  I	  �	  �	  
  <
  t
  �
  �
  %  ^  �  �    ?  x  �  �    V  �  �    H  �  �  �  2  j  �  �  �  �  )  H  u  �  �    H  �  �  �  �  8  s  �  �    R  �  �    E  |  �  �  #  Y  �  �  �  2	  e	  �	  �	  
  @
  n
  �
  �
    K  ~  �  �  &  ]  �  �  �  1  i  �  �    ;  s  �  �  �  �  �    K  p  �  �  �    C  q  �  �  �  7  x  �  �  !  X  �  �    =  p  �  �     '  a  �  �  �  "	  F	  �	  �	  �	  
  K
  z
  �
  �
    ;  j  �  �    F  t  �  �    F  v  �  �    X  x  �  �  C  H  m  �  �  �  �  5  q  �  �  �  2  g  �  �  �  2  `  �  �  �    F  u  �  �  �  !  V  �  �  �  	  E	  z	  �	  �	  
  :
  t
  �
  �
  	  6  m  �  �  
  >  s  �  �  
  ?  a  [  q  �  �  �  �    N  x  �  �  �    B  w  �  �  �  $  I  ~  �  �    *  H  �  �    +  M  s  �  �  %  X    �  �  	  L	  �	  �	  �	  
  @
  }
  �
  �
    <  q  �  �    :  g  �  @  M  _  j  i  q  t  �  �  �  "  F  a  �  �  �  �  /  u  �  �  �     =  �  �  �    ,  c  �  �     =  _  �  �     K  m  �  �  	  O	  ~	  �	  �	  �	  C
  �
  �
  �
  �
  5  y  �  �    %      2  ,      <  C  h  p  �  �  �    ]  �  �  �  �  4  �  �  �  �    i  �  �  �    Q  �  �    ,  I  �  �  $  N  a  �  �  	  X	  �	  �	  �	  
  Q
  �
  �
  �
  �
  =  �  �  �  �  �  �  �  �  �  �  �  �  �  "  �  �  |  �    L  �  �  �  �  I  �  �  �  �  #  |  �  �  �    Y  �  �    )  H  �  �    M  \  �  �  	  P	  }	  �	  �	  
  O
  �
  �
  �
  �
  >  �  �  �  n  /  �  �  X  J  k  ]  �  �  k  t  g  �  
  _  �  �  �  �  Q  �  �  �  �  D  �  �  �    B  �  �    *  O  �  �    D  d  �  �  	  U	  |	  �	  �	  
  \
  �
  �
  �
    ]  �  �  �    ,  ,  �  �  �  �  �  �  �  V  �  �  �  �  +  u  �  �  �    f  �  �  �    [  �  �  �    X  �  �    5  _  �  �  (  O  q  �  �  -	  a	  �	  �	  �	  /
  n
  �
  �
  �
  0  s  �  �    7  D  ,  \  �    V  C  U  t  �  �  �  �  9  �  �  �  �  &  l  �  �  �  !  Z  �  �    .  W  �  �    ;  a  �  �  "  P  u  �  �  %	  _	  �	  �	  �	  #
  e
  �
  �
  �
  (  j  �  �  �  0  m  ,  ,  j  �  .  m  ]  �  �  �  0  c  �  �  �    3  ]  �  �  �     M  |  �  �  !  D  p  �  �  &  O  w  �  �  #  Y  �  �  �  	  ]	  �	  �	  �	  
  a
  �
  �
  �
  &  e  �  �    2  k  �  f  �  �  �  M  j  }  �  �  ?    �  �  �  '  n  �  �  �    [  �  �  �    M  �  �  �    D    �  �    >  v  �  �  	  :	  o	  �	  �	  
  A
  s
  �
  �
    F  y  �  �    M    �  �    �      T  m  �    C  i  �  �    Z  �  �  �  %  f  �  �    =  t  �  �  '  U  �  �  �  2  a  �  �  	  <	  g	  �	  �	  �	  7
  h
  �
  �
  �
  1  f  �  �  �  ,  c  �  �  �  .  d  �  r  7  /  O  m  �  �  3  d  �  �    Y  �  �  �  >  ~  �  �  $  h  �  �    N  �  �  �  6  q  �  �  	  _	  �	  �	  �	  /
  e
  �
  �
    >  r  �  �    ?  q  �  �  
  .  _  �  �  �  3  `  a  ]  p  �  �    F  �  �    C  �  �    :  t  �  �  -  f  �  �    Z  �  �    Q  �  �  	  E	  �	  �	  �	  7
  t
  �
  �
  (  e  �  �    S  �  �    >  s  �  �    <  q  �  �  �  f  a  p  �  +  8  d  �  �    3  j  �  �  "  W  �  �    O  �  �    R  �  �    V  �  �  	  Q	  �	  �	  

  I
  �
  �
    F  �  �    A  �  �  �  9  v  �  �  .  j  �  �    a  �  �  Z  �  �    ;  r  �  �  "  S  �  �  �  6  n  �  �     \  �  �    Q  �  �    E  �  �  �  :	  {	  �	  �	  4
  w
  �
  �
  0  q  �  �  .  l  �  �  ,  h  �  �  '  d  �  �     ^  �  �    ^  �    A  l  �  �    X  �  �  �  F    �  �  -  q  �  �    Z  �  �    I  �  �  	  B	  ~	  �	  
  ;
  v
  �
  �
  4  o  �  �  *  h  �  �     `  �  �    W  �  �    N  �  �  	  G  c  �  P  r  �  �  
  0  s  �  �  
  e  �  �    L  �  �    M  �  �    G  �  �  	  D	  }	  �	  �	  @
  |
  �
  �
  :  y  �  �  0  r  �  �  (  g  �  �     ^  �  �    W  �  �    O  �  �  �  �  �  �  �  )  c  �  �    S  �  �  �  "  P  �  �    8  t  �    6  j  �  �  6	  n	  �	  �	  .
  l
  �
  �
    Z  �  �    B  �  �  �  2  m  �  �  #  _  �  �    R  �  �    A  �  �  �  *  �  �  &  �  �  �  	  Z  �  �  �  @  �  �  �  0  b  �  �    K  �  �  �  +	  ^	  �	  �	  	
  B
  x
  �
  �
  #  _  �  �    B    �  �  +  f  �  �    S  �  �    P  �  �    �  �  �    �  d  �  �    �  �  a  �  �  �  )  x  �  �  $  V  �  �    M  {  �  �  6	  l	  �	  �	  
  O
  �
  �
  �
  .  i  �  �    H  �  �  �  *  d  �  �    H  �  �  �  0  h  �  �  �  �  �  m  �  �  �  �  '  �  �  �  �  '  d  �  �  �  +  [  �  �  �  1  b  �  �  	  >	  t	  �	  �	  
  M
  �
  �
  �
  "  ^  �  �    7  q  �  �    N  �  �  �  0  f  �  �    H    �  �  �    �  �  �  �    �  �  �    3  �  �    ,  Y  �  �    D  o  �  �  &	  W	  �	  �	  �	  1
  g
  �
  �
    @  w  �  �    R  �  �  �    U  �  �  �  "  Z  �  �  �  *  a  �  �    �  �  O  �  �  �  C  �  �  �  �  b  �  �    /  y  �    =  d  �  �  /	  a	  �	  �	  
  N
  �
  �
  �
  *  j  �  �    J  �  �  �  0  j  �  �    M  �  �  �  6  k  �  �    I  �  �  �  {  �  �  �  �  �  h  �  �  �    {  �  �  )  e  �  �    T  �  �  	  J	  ~	  �	  �	  8
  k
  �
  �
    W  �  �  �  :  u  �  �     [  �  �    @  }  �  �  *  b  �  �    J  �  �  �  5  Z  j  ~  �  �  �  @  �  �  �  =  �  �  �  !  f  �  �    N  �  �  �  .	  g	  �	  �	  
  Q
  �
  �
  �
  *  f  �  �    Q  �  �  �  1  j  �  �    M  �  �  �  3  k  �  �  .  h  �  �      |  �  �  �    m  �  �    E  x  �  �  ,  _  �  �    J    �  �  1	  p	  �	  �	  
  W
  �
  �
    @  �  �  �  2  m  �  �  (  ^  �  �    N  �  �  �  8  q  �  �    Y  �  �    D    I  |  �  �  	  2  {  �  �  ,  a  �  �    P  �  �    >  r  �  �  "	  ]	  �	  �	  �	  ?
  }
  �
  �
    [  �  �    =  z  �  �  )  _  �  �    K  �  �  �  5  m  �  �    V  �  �  �    �  4  �  �  	  %  H  �  �  !  A  h  �  �  2  \  �  �    @  q  �  �  	  P	  �	  �	  �	  "
  c
  �
  �
     9  y  �  �    T  �  �    ;  q  �  �  %  [  �  �    D  |  �  �  '  d  �  �  �  ,  �  �  �  
  @  �  �  �     K  �  �    ;  g  �  �  )  ^  �  �  	  P	  �	  �	  �	  ;
  {
  �
  �
  (  k  �  �    U  �  �    M  �  �    B  ~  �  �  6  r  �  �  )  g  �  �    �  �  %    |  �  �    K  �  �    8  �  �    B  n  �    D  z  �  �  A	  }	  �	  �	  8
  {
  �
  �
  /  s  �  �  -  m  �  �  )  f  �  �  &  a  �  �    \  �  �    S  �  �    F  �  �  �    (  h  �  �  �  J  �  �    :  �  �    L  �  �    S  �  �  	  W	  �	  �	  
  S
  �
  �
    Q  �  �    K  �  �    C  �  �  �  <  z  �  �  1  m  �  �    X  �  �    N  R  U  �  �  �  L  �  �  �  *  z  �     3  v  �    8  s  �  �  >  u  �  �  7	  t	  �	  �	  4
  t
  �
  �
  +  j  �  �    V  �  �    I  �  �  �  4  l  �  �    U  �  �    B  w  �  �  �  O  �  �  �  +  t  �  �    P  �  �  
  ?  �  �    =  w  �  �  5  m  �  �  $	  c	  �	  �	  
  P
  �
  �
  �
  +  e  �  �    L  �  �  �  &  \  �  �  
  ?  t  �  �    S  �  �  �  �  �  L  o  �  �  �  ,  n  �  �    Y  �  �    >  |  �  �  ,  d  �  �    L  w  �  �  	  F	  r	  �	  �	  
  K
  {
  �
  �
    J  {  �  �    Q  �  �  �    S  �  �  �  $  \  �  �  �  �  �    P  v  �  �  �  :  r  �  �  �  ?  z  �  �    M  �  �  �    K  �  �  �    ?  x  �  �  �  ,	  k	  �	  �	  �	  $
  ]
  �
  �
  �
  .  b  �  �    6  i  �  �    9  h  �  �    <  <  <  �    6  p  �  �  �    `  �  �  �    <  d  �  �    <  Z  �  �  �  2  W  �  �  �    F  {  �  �  �  	  K	  	  �	  �	  
  >
  q
  �
  �
  �
  $  Z  �  �  �  &  U  �  �  �  $  K  �  �  �  �  �  :  p  ~  �  �      I    �  �  �    R  x  �  �  �  /  R  v  �  �    4  X  x  �  �    7  `  �  �  �  	  R	  �	  �	  �	  
  A
  y
  �
  �
  �
  /  f  �  �    6  d  �  �  	  �  �  �  �    '  Y  �  �  �  �  �  !  K  V  �  �  �  �    9  q  �  �      (  ^  �  �    0  O  }  �    <  `  |  �  �  0	  d	  �	  �	  �	   
  c
  �
  �
  �
    N  �  �  �    A  �  �  �  �  �  {  �    6  5  A  I  v  �  �  �  �  �  %  e  �  �  �  �  &  s  �  �  �    Q  �  �    +  J  �  �    ?  ]    �  	  G	  q	  �	  �	  �	  >
  {
  �
  �
  �
  /  t  �  �  �  !  7  M  a  �  �  v  �  �  �  �  �  �  �  $  O  �  �  �  �  C  �  �  �  �  !  y  �  �  �    _  �  �    -  S  �  �  %  M  a  �  �  $	  X	  ~	  �	  �	  
  V
  �
  �
  �
  �
  ?  �  �  �  �       '  O  ;  �  _  �  �  �  �  �  �    L  �  �  �  �  ;  �  �  �  �  &  t  �  �  �  $  [  �  �    0  X  �  �  $  L  d  �  �  	  W	  ~	  �	  �	  
  K
  �
  �
  �
  �
  :  �  �  �    �  }    /  +  L  G  v  �          >  �  �  �  �    `  �  �  �    K  �  �    !  H  �  �    9  Z  �  �    G  n  �  �  	  N	  	  �	  �	  
  N
  �
  �
  �
    P  �  �  �    S  g  k  �  3  p  �  �  �  �  L  x  z  �  �  �  '  6  c  �  �  
  4  Q  {  �  �  -  O  t  �  �  '  X  }  �  �    Y  �  �  �  	  V	  �	  �	  �	  
  U
  �
  �
  �
    R  �  �  �  #  X  �  }  �    @  �  �  �  �  5  u  �  �  �    Y  �  �  �    C  y  �  �  �  *  d  �  �  �    P  �  �  �  
  E  �  �  �  	  ?	  {	  �	  �	  
  =
  o
  �
  �
    9  n  �  �    F  v  �  �  %    0  }  �  �  �    [  �  �  �    W  �  �  �    I  �  �  �    G  �  �  �    >  t  �  �    ?  p  �  �  	  ;	  i	  �	  �	  
  :
  f
  �
  �
    B  n  �  �    E  t  �  �    G  $  I  k  �  �  �  E  f  �  �  �    W  �  �  �    I  �  �  �  $  L  �  �  �  -  V  �  �  �  .  \  �  �  �  ,	  _	  �	  �	  �	  '
  ^
  �
  �
  �
  )  b  �  �  �  ,  d  �  �  �  /  f  �  b  t  �  �  �  .  n  �  �  �  H  �  �  �    R  �  �     2  n  �  �    J    �  �  (  `  �  �  �  4	  l	  �	  �	  
  L
  �
  �
  �
  "  P  �  �  �     N  |  �  �    P  �  �  �    S  �  �  �  �  0  m  �  �  �  F  �  �  �  $  h  �  �    M  �  �    >  u  �  �  *  _  �  �  	  F	  }	  �	  �	  5
  l
  �
  �
    X  �  �  �  .  c  �  �  �  ,  b  �  �  �    O  �  �  �  �  �  �  >  l  �  �  �  D  �  �  �  +  r  �  �    X  �  �    I  �  �    C  {  �  �  7	  r	  �	  �	  '
  e
  �
  �
    U  �  �    D  �  �  �  4  p  �  �  "  Z  �  �  �  '  V  �  �  �  �    V  �  �  �  1  z  �  �    b  �  �  	  S  �  �     I  �  �  �  C  �  �  �  @	  �	  �	  �	  9
  y
  �
  �
  5  v  �  �  .  o  �  �  '  e  �  �    [  �  �    O  �  �    I  �    X  `  f  �  �  "  k  �  �    K  �  �    7  �  �  �  /  n  �  �  -  g  �  �  *	  b	  �	  �	  $
  ]
  �
  �
  !  ]  �  �    Z  �  �    U  �  �    N  �  �    G  �  �    ?  ~  �    b  �  �  �    /  y  �  �    m  �  �    Q  �  �  #  P  �  �    S  �  �  	  P	  �	  �	  
  H
  �
  �
  �
  ;  |  �  �  1  s  �  �  )  h  �  �  !  ^  �  �    S  �  �  
  G  �  �  0  b  �  �  �  P  �  �  �  3  P  t  �  �  '  X  �  �    M  �  �    L  �  �  	  E	  }	  �	  �	  :
  w
  �
  �
  /  m  �  �  !  b  �  �    R  �  �    @  {  �  �  /  j  �  �  #  d  �  �  �  �  �    i  �  �  
  F  z  �  �  ;  f  �  �    7  r  �  �    L  �  �  �  1	  g	  �	  �	  
  Q
  �
  �
  �
  5  q  �  �    Y  �  �    C    �  �  1  m  �  �     [  �  �    H  �    *  �  B  }  �  �    P  �  �  	  D  |  �  �  =  t  �  �    N  �  �  �  /	  e	  �	  �	  
  J
  �
  �
  �
  *  e  �  �    L  �  �  �  )  _  �  �  	  >  r  �  �    T  �  �  �  2  �  4  t  �  �  �    &  _  t  �  �  !  M  �  �  �  4  j  �  �    Y  �  �  �  7	  s	  �	  �	  
  R
  �
  �
  �
  4  n  �  �    O  �  �  �  4  m  �  �    O  �  �  �  3  j  �  �    L  Z  I  k  �    &  M  �  �    (  J  z  �  �    <  u  �  �    A  t  �  �  	  J	  �	  �	  �	  "
  Y
  �
  �
  �
  4  k  �  �    G    �  �  &  \  �  �    ;  s  �  �    R  �  �  �  1  D  �  �  �    `  �  �    =  s  �  �    N  �  �  �    T  �  �  �  (	  ]	  �	  �	   
  5
  i
  �
  �
    B  w  �  �    Q  �  �  �  !  V  �  �  �  *  ]  �  �  �  3  g  �  �    =  r  =  T  �  (  Y  �  �  �  #  \  �  �    9  d  �  �    P  �  �  �  2	  k	  �	  �	  
  M
  �
  �
  �
  '  f  �  �    D  �  �  �  +  b  �  �    I  ~  �  �  .  e  �  �    H  �  �  �  (  �  �  �  �  7  W  �  �    .  Z  �  �  0  `  �  �    S  �  �  	  B	  u	  �	  �	  "
  ^
  �
  �
    @  z  �  �  #  ^  �  �    D  ~  �  �  +  d  �  �    L  �  �  �  2  l  �  �    U  ~  �  �  �    $  �  �  �  .  d  �  �    U  �  �    ;  q  �  �  	  N	  �	  �	  �	  9
  q
  �
  �
    L  �  �    8  q  �  �    S  �  �  �  8  p  �  �    U  �  �    L  �  �  �  3  �  �  4  �  �  �  �  0  {  �  �    L  �  �    <  n  �  �  2	  b	  �	  �	  
  W
  �
  �
  �
  >  {  �  �    Z  �  �    ;  {  �  �  '  ^  �  �    I    �  �  3  j  �  �    U  �  �  �  �    S  �  �  �  )  w  �  �    I  �  �    3  h  �  �  "	  S	  �	  �	  

  C
  u
  �
  �
  '  c  �  �    B  �  �  �     ^  �  �  
  ?  {  �  �  *  _  �  �    J    �  �  1  j  �  �  �  �  K  �  �  �    P  �  �  �  %  b  �  �    @  s  �  �  (	  W	  �	  �	  �	  8
  m
  �
  �
    K  �  �  �  #  _  �  �    :  t  �  �    R  �  �  �  6  l  �  �    Q  �  �  �  3  �  �  �  <  �  �  �  �  @  p  �  �    H  y  �  �  *  [  �  �  	  =	  s	  �	  �	  
  Y
  �
  �
    >  y  �  �  %  a  �  �    I  �  �  �  4  n  �  �  !  Z  �  �    F    �  �  /  j  �  �  �    4  i  �  �    >  �  �  �  %  Z  �  �    D  {  �  �  1	  o	  �	  �	  "
  \
  �
  �
    N  �  �    =  {  �  �  -  i  �  �    U  �  �    @  x  �  �  )  a  �  �    F  ~  q  �  �  �    [  �  �  �     T  �  �    <  x  �  �  5  q  �  �  %	  _	  �	  �	  
  U
  �
  �
  	  F  �  �  �  0  l  �  �    J  �  �  �  /  j  �  �    J  �  �  �  %  \  �  �  �  �      �  �  �    Q  �  �  �  /  i  �  �    T  �  �  �  =  z  �  �  /	  j	  �	  �	  
  Y
  �
  �
  �
  7  p  �  �    8  j  �  �    M  �  �  �  #  V  �  �  �  9  o  �  �  �          i  �  �  �  �    P  �  �  �  3  i  �  �    F  {  �  �    Y  �  �  	  :	  f	  �	  �	  
  6
  a
  �
  �
  �
  '  Z  �  �    9  n  �  �  �  2  i  �  �  �  4  j  �  �  �  #  J  P  P  �  &  Y  l  �  �  �    F  z  �  �    C  x  �  �    @  �  �  �    =  l  �  �  �  	  K	  �	  �	  �	  

  <
  p
  �
  �
    2  c  �  �  �  2  d  �  �  �  .  c  �  �  �  +  _  �  �  �  �  �      9  x  �  �  �    H  w  �  �  �  $  V  �  �  �  
  <  k  �  �  �     U  z  �  �  �  :	  s	  �	  �	  �	  )
  d
  �
  �
  �
  '  X  �  �     0  \  �  �  �    S  �  �  �  �  �  �  �  �  �  �    C  i  �  �  �    "  ;  _  �  �    *  D  i  �  �    =  `  �  �  �  ,  \  �  �  �  �  &	  Y	  �	  �	  �	  
  E
  {
  �
  �
  �
  )  ]  �  �  �     R  �  �  �    J  x  �  �  �  �  �  �  �  �    /  S  �  �  �  �    L  �  �  �  �  '  D  h  �  �  �    >  \  q  �  �    E  h  �  �  �  6	  g	  �	  �	  �	  "
  ^
  �
  �
  �
    K  �  �  �    B  {  �  �  k  j  a  Y  n  {  �  �  �  �  �    ]  r  �  �  �  �  �    ?  m  �  �  �      H  �  �    !  ;  m  �  �  2  P  k  �  �  *	  \	  	  �	  �	  
  ]
  �
  �
  �
    I  �  �  �    ;  }  J  F    �  �    )  [  �  �  �  �  �  �  �  �     0  k  �  �  �  �  8  �  �  �  �  &  m  �  �    2  ^  �  �  +  M  g  �  �  %	  \	  	  �	  �	  
  Z
  �
  �
  �
    J  �  �  �    :  '  "  �  �  �  �  �  F  j  _  �  �  �  �  �  �    �  C  �  �  �  �  '  r  �  �    $  Z  �  �    0  S  �  �    K  ^  �  �  	  O	  y	  �	  �	  �	  >
  ~
  �
  �
  �
  &  p  �  �  �    �    �  �  �  �  �    O  e  �  �  �    6  @  N  P  �  �  
  .  ;  `  �  �    ;  [  �  �    C  b  �  �    K  x  �  �  �  >	  	  �	  �	  �	  4
  w
  �
  �
    4  n  �  �    >  m  f  �  $  �  �  �  �  &  l  �  �  �  �     k  �  �  �  �  )  a  �  �  �     <  r  �  �  �  &  n  �  �  �  "  _  �  �  �  	  S	  �	  �	  �	  
  O
  �
  �
  �
    N  �  �  �  )  U  �  �  k  �  �  .  6  &  ,  T  �  �  �    =  {  �  �  �  '  `  �  �  �  !  N  �  �  �    >  r  �  �  
  0  ]  �  �  	  -	  Z	  �	  �	  �	  *
  V
  �
  �
  �
  +  X  �  �  �  "  S  �  �  �  %  y  �  �  @  }  �  �  �  �    0  L  �  �    -  S  �  �  �  +  M  v  �  �     P  y  �  �    D  o  �  �  	  A	  p	  �	  �	  
  :
  m
  �
  �
  �
  +  a  �  �  �  $  _  �  �  �  '  ]  �  �  �  �  7  �  �  �  �  6  m  �  �  �    I  x  �  �  
  >  m  �  �    8  l  �  �  �  ,  i  �  �  �  )	  b	  �	  �	  �	  %
  [
  �
  �
  �
  "  V  �  �  �  )  Z  �  �  �  -  \  �  �  �  �  �  .  N  ~  �  �    T  �  �  �    S  �  �  �    M  �  �  �  !  O  �  �  �  !  P  �  �  �  	  N	  ~	  �	  �	  
  L
  |
  �
  �
    J  }  �  �    Q  �  �  �  !  V  �  �  �  %  Z    ,  `  z  �  �  (  U  �  �     <  v  �  �    V  �  �  �  5  n  �  �    J  �  �  �  &	  _	  �	  �	  �	  1
  m
  �
  �
    ;  r  �  �    7  m  �  �    2  j  �  �    6  k  �  �  	  �  v  p  �  �  #  U  �  �  �  =  r  �  �  #  e  �  �    K  �  �  �  7  s  �  �  !	  Z	  �	  �	  

  A
  
  �
  �
  1  i  �  �    H  {  �  �    I  {  �  �    J  u  �  �    8  m  �  �  �  �  �  
  Q  p  �  �  1  n  �  �    a  �  �    M  �  �    <  z  �  �  4	  o	  �	  �	  +
  e
  �
  �
    Z  �  �    L  �  �  �  <  y  �  �  *  f  �  �    >  p  �  �    4  f  �  �  �  �  K  t  �  �    Z  �  �  
  I  z  �    ?  s  �  �  8  o  �  �  6	  m	  �	  �	  /
  j
  �
  �
  '  g  �  �    ]  �  �    S  �  �    J  �  �    A    �  �  9  t  �  �  2  �  �  �    �  �  �  �  O  �  �  �  ,  b  �  �    P  �  �    N  �  �  		  F	  }	  �	  �	  ;
  w
  �
  �
  /  n  �  �  #  b  �  �    R  �  �  
  E  �  �  �  8  t  �  �  +  i  �  �    �    T  �  �  �  �    m  �  �    K  �  �    :  u  �  �  %  [  �  �  		  D	  {	  �	  �	  -
  h
  �
  �
    U  �  �    =  z  �  �  %  `  �  �    K  �  �  �  8  r  �  �  (  g  �  �  �  �  v  �  �  �  9  U  �  �      K  �  �    @  w  �  �  8  j  �  �  	  V	  �	  �	  �	  5
  n
  �
  �
    M  �  �  �  -  h  �  �    J  �  �  �  1  i  �  �    Q  �  �    ?  x  �  �  �  �  �  �  �  )  �  �       ]  �  �    E  u  �  �  %  \  �  �  �  3	  l	  �	  �	  
  D
  
  �
  �
    W  �  �  �  4  l  �  �    K  �  �  �  .  e  �  �    G  ~  �  �  )  a  �  �  �  �  
  �    g  �  �  	  4  r  �    2  [  �  �    V  �  �  �  5	  o	  �	  �	  
  B
  y
  �
  �
    R  �  �  �  0  f  �  �    D  z  �  �  "  Y  �  �  �  7  o  �  �    P  �  �  �  �    P  �  �  �  �    %  F  �  �     :  a  �  �  1  \  �  �  	  H	  |	  �	  �	  
  ]
  �
  �
  �
  2  o  �  �    J  �  �  �  +  a  �  �    A  w  �  �    V  �  �  �  6  n  �  �  �  �    �  �  �  
  &  s  �  �    8  a  �  �  �  :  f  �  �  �  2	  l	  �	  �	  �	  7
  v
  �
  �
    A  �  �  �    P  �  �  �  0  c  �  �    E  w  �  �  "  Y  �  �  �  3  l  �  �  �    N  �  �  �    P  �  �  	  %  Z  �  �  !  C  l  �  �  *	  X	  �	  �	  �	  0
  f
  �
  �
  �
  8  q  �  �  
  D  }  �  �    S  �  �  �  $  [  �  �  �  .  d  �  �    9  o  �  �    �  �  B  �  �  �    C  �  �    4  d  �  �  $  T  �  �  	  B	  t	  �	  �	  #
  _
  �
  �
  �
  <  y  �  �    V  �  �  �  5  q  �  �    R  �  �    9  n  �  �    U  �  �  �  9  q  �  �  �    x  �  �    J  �  �    =  w  �  �  -  _  �  �  	  P	  �	  �	  �	  2
  l
  �
  �
  
  M  �  �  �  (  j  �  �    G  �  �  �  1  h  �  �     T  �  �    @  v  �  �  $  `  �  �  �  �  1  �  �  �    C  �  �  �  *  Y  �  �    I  u  �  �  0	  a	  �	  �	  
  I
  ~
  �
  �
    ]  �  �  �  @  }  �  �  #  [  �  �    A  y  �  �  *  a  �  �    L  �  �  �  9  t  �    >  v  �  �    Q  ~  �  �  7  n  �  �    T  �  �  �  9	  u	  �	  �	  
  [
  �
  �
    =  �  �  �  +  `  �  �    N  �  �  �  ;  q  �  �    Z  �  �     <  x  �  �    [  �  �    �  /  \  �  �    H  w  �  �  -  i  �  �    M  �  �  �  3	  l	  �	  �	  
  O
  �
  �
  �
  0  m  �  �    M  �  �  �  6  l  �  �    U  �  �    <  t  �  �    Z  �  �    =  x  �  �  �    =  �  �    8  ^  �  �    P  z  �  �  -  e  �  �  �  :	  t	  �	  �	  
  H
  �
  �
  �
  !  [  �  �    8  p  �  �    O  �  �  �  2  g  �  �    H    �  �  &  _  �  �    =  v  �    6  �  �  �  #  H  �  �  �  0  ^  �  �    A  t  �  �  	  W	  �	  �	  �	  4
  p
  �
  �
    N  �  �  �  .  i  �  �    K  �  �  �  /  g  �  �    K  �  �  �  .  e  �  �    G  }  �  	  "  ^  �  �     0  _  �  �    =  l  �  �  *  V  �  �  	  E	  w	  �	  �	  #
  _
  �
  �
    A  {  �  �  "  [  �  �     :  v  �  �    R  �  �  �  /  g  �  �    B  z  �  �      �  �    5  _  �  �    0  p  �  �    O  �  �    7  s  �  �  	  P	  �	  �	  �	  .
  a
  �
  �
    ?  v  �  �    Q  �  �  �  $  b  �  �  �  5  m  �  �  	  @  u  �  �    =  ?  A  A  {  �  �    G  x  �  �  	  C  ~  �  �  !  P  �  �  �  !  Z  �  �  �  %	  a	  �	  �	  �	  +
  a
  �
  �
    2  ]  �  �     /  c  �  �    9  j  �  �    7  k  �  �    7  k  }  �  �  �  m  �  �  �  �  7  �  �  �    -  l  �  �  �  -  ]  �  �  �     V  �  �  �  	  K	  |	  �	  �	  
  4
  Z
  �
  �
  �
    L  �  �  �  )  Q  �  �  �    P  �  �  �    L    �  �  �  �  �  :  t  �  �  �  �  5  S  �  �  �    9  ]  �  �  �    >  }  �  �  �  (  Z  �  �  �  �  *	  `	  �	  �	  �	  
  @
  s
  �
  �
    3  e  �  �    0  Y  �  �  �  -  ^  �  �  �  &  \  a  a    F  l  }  �  �  �  �  )  R  �  �  �  �    5  Y  {  �  �    5  [  t  �  �    ;  a  �  �  �  	  W	  �	  �	  �	  
  D
  
  �
  �
    5  t  �  �  
  3  f  �  �  �  &  Y  �  �  �  �  �      3  e  �  �  �  �  �    1  ;  L  m  �  �  �  "  ;  \  �  �    ,  K  w  �  �    B  l  �  �  �  	  A	  n	  �	  �	  �	  &
  `
  �
  �
  �
  
  A  y  �  �    4  k  �  �  �  -  [  �  �  �  �    E  N  W  Z  t  �  �  �  �      R  �  �  �    %  E  f  �  �  �    0  L  [  �  �    ;  X  }  �  �  1	  `	  �	  �	  �	  
  \
  �
  �
  �
  
  K  �  �  �    ?  |  �  �  �  �  �  �  �  �  �  �      %  \  �  �  �  �      (  ?  \  z  �  �        Y  �  �    '  K  �  �    A  Z    �  	  F	  p	  �	  �	  �	  :
  w
  �
  �
  �
  )  k  �  �  �    Y  �  �  �  �  �  �  �  �  �  �      J  o  �  �  �  �  �      )  3  K  �  �    #  @  x  �    -  H  n  �  �  0  [  y  �  �  '	  f	  �	  �	  �	  
  ]
  �
  �
  �
    K  �  �  �    B  �  y  ~  }  �  �  �  �  �  �  �  �  �  J  {  �  �  �  �  '  ^  t  �  �  �    N  k    �  �  +  c  �  �  �    Q  �  �  �  �  9	  y	  �	  �	  �	  $
  f
  �
  �
  �
    R  �  �       G  �    y  ~  g  �  �  �        "  )  V  �  �  �      \  �  �  �  �    W  �  �  �    9  u  �  �  �  $  ^  �  �  	  .	  b	  �	  �	  
  .
  [
  �
  �
    2  ]  �  �  �  3  `  �  �     �  7  �    �  �  �  �  N  ]  n  q  �  �    :  W  v  �  �    A  a  �  �  �  /  W    �  �  +  U  }  �  �  	  I	  s	  �	  �	  
  A
  o
  �
  �
    9  j  �  �  �  1  g  �  �  �  '  ]  �  6  �  �  �  �  �    b  �  �  �    >  b  �  �  �    K  ~  �  �    =  s  �  �  �  -  f  �  �  �  	  V	  �	  �	  �	  
  O
  �
  �
  �
    D  |  �  �    ?  r  �  �    6  i  �  �  �  E  �  �  �    B  {  �  �  �    Q  �  �  �    H  ~  �  �    7  k  �  �    1  f  �  �  �  #	  T	  �	  �	  �	  &
  T
  �
  �
  �
  $  S  �  �  �    I  x  �  �    O    �  �    J  Z  q  �  �  �    W  �  �    0  _  �  �    *  O  �  �  �  +  R  �  �  �  '  P  }  �  �  #	  T	  �	  �	  �	  
  P
  ~
  �
  �
    L  }  �  �    G    �  �    J  �  �  �    K  �  �  k  �  �  �     l  �  �  �  "  U  �  �     2  ]  �  �  �  3  d  �  �  �  4  h  �  �  �  2	  i	  �	  �	  �	  /
  f
  �
  �
  �
  ,  c  �  �  �  -  g  �  �    3  h  �  �  
  ;  m  �  �    �  �  �     R  �  �  �  4  e  �  �    K  �  �    7  h  �  �    L  �  �  �  -	  b	  �	  �	  
  ;
  o
  �
  �
    S  �  �  �  %  X  �  �  �  "  V  �  �  �    S  �  �  �     V  �  �  #  �  �  ;  �  �  �    ]  �  �    N  �  �    E  y  �  �  1  n  �  �  	  V	  �	  �	  
  <
  w
  �
  �
  &  e  �  �    L  �  �  �  .  a  �  �  �  ,  _  �  �  �  &  M  �  �  �    Q    �  '  g  �  �    A  �  �    =  u  �  �  7  k  �  �  ,  c  �  �  	  Z	  �	  �	  
  L
  �
  �
    >  ~  �  �  2  o  �  �  '  b  �  �    U  �  �  	  E    �  �    T  �  �  �      S  t  �  �  �  7  l  �  �    V  �  �    H  y  �  �  ;  t  �  �  +	  i	  �	  �	  
  ^
  �
  �
    N  �  �    @  �  �  �  4  s  �  �  )  f  �  �    X  �  �    H  �  �  �  5  s  �  n  w  �    .  T  �  �    I  �  �  �    X  �  �    ?  w  �  �  '	  c	  �	  �	  
  N
  �
  �
  �
  6  t  �  �     \  �  �    F  �  �  �  4  n  �  �     Z  �  �    G  �  �  �  5  q  �  �  !  C  X  m  �  �  4  d  �  �    R  �  �  �  3  p  �  �  	  J	  �	  �	  �	  (
  a
  �
  �
    A  |  �  �  #  ]  �  �  
  B  |  �  �  *  _  �  �    E  |  �  �  (  b  �  �    t  �  �  .  F  �  �  �  0  \  �  �  �  '  c  �  �    A  �  �  �  &	  `	  �	  �	  
  B
  {
  �
  �
  %  ]  �  �    >  w  �  �  "  Z  �  �    >  s  �  �    U  �  �  �  2  k  �  �    2  f  C  ?  q  �  �  (  b  �  �  �  ;  u  �  �    D  s  �  �  	  K	  �	  �	  �	  %
  Z
  �
  �
    9  n  �  �    N  �  �  �  +  c  �  �  	  A  z  �  �  !  Y  �  �     8  p  �  �    A  y  �  �  �  �    F  l  �  �    X  �  �  �  6  |  �  �  	  S	  �	  �	  �	  .
  e
  �
  �
    F  {  �  �  $  [  �  �    9  q  �  �    F  |  �  �    T  �  �  �  -  c  �  �    ;  N  �  �  �     ,  �  �  �  �  �  ;  }  �  �  
  D  �  �  �  "	  ]	  �	  �	  	
  =
  w
  �
  �
  #  W  �  �    ;  q  �  �    R  �  �  �  0  i  �  �    F  |  �  �  !  Z  �  �    7  o  �  �  �  �    Z  �  �  �  0  ^  �  �  �  $  M  �  �  �  #	  Q	  �	  �	  �	  )
  Y
  �
  �
    9  i  �  �    H  {  �  �    X  �  �  �  /  i  �  �    B  {  �  �     V  �  �  �  4  j  �  W  �  �  1  5  f  �  �  *  W  {  �  �  5  l  �  �  �  @	  {	  �	  �	  
  K
  �
  �
  �
  !  Y  �  �    4  j  �  �    H  }  �  �  "  V  �  �  �  1  d  �  �    >  s  �  �    L  �  L  R    �  �  (  `  �  �     R  �  �  �  5  p  �  �  
	  N	  �	  �	  �	  )
  h
  �
  �
    F  �  �  �  /  b  �  �    L    �  �  2  i  �  �    L  �  �  �  +  f  �  �    E  �  �  �  3  9  _  �    @  f  �  �     W  �  �  �  ?  z  �  �  	  ^	  �	  �	  �	  6
  x
  �
  �
    Q  �  �    :  p  �  �  )  [  �  �    H  |  �  �  *  i  �  �    J  �  �  �  -  i  �  �      3  s  �    @  ]  �  �    K  z  �  �  &  g  �  �  �  7	  x	  �	  �	  
  N
  �
  �
  �
  -  f  �  �    H  �  �  �  7  k  �  �    S  �  �  �  5  p  �  �    R  �  �    A  |  �  �  �  �    V  {  �    .  b  �  �    G  {  �  �  +	  `	  �	  �	  
  ?
  v
  �
  �
    Z  �  �    <  y  �  �  $  ^  �  �    E    �  �  .  g  �  �    Q  �  �  �  9  q  �  �    U  �  �  �  
  6  q  �  �    O  �  �     6  k  �  �  	  T	  �	  �	  
  =
  t
  �
  �
    Y  �  �     9  t  �  �    U  �  �    :  r  �  �    W  �  �    =  u  �  �  !  [  �  �    ?  y  �  �    ,  [  �  �    <  m  �  �    M  �  �  �  '	  [	  �	  �	  �	  1
  g
  �
  �
    >  w  �  �    M  �  �  �  %  \  �  �    5  k  �  �    F  {  �  �  !  V  �  �  �  1  f  �  �  �  �  �    7  t  �  �    C  y  �  �    H  w  �  �  	  T	  �	  �	  �	  "
  ^
  �
  �
  �
  .  f  �  �    9  p  �  �    J  �  �  �    X  �  �  �  0  g  �  �    @  v  �  �    D  E  t  �  �  �    D  t  �  �    0  k  �  �    B  q  �  �  	  :	  s	  �	  �	  
  ?
  x
  �
  �
    N  �  �  �  '  Y  �  �  �  /  h  �  �    >  v  �  �    H  ~  �  �    O  �  �  �  �  @  c  �  �  �    <  k  �  �    ,  T  �  �  �  "  S  �  �  �  	  X	  �	  �	  �	  "
  T
  �
  �
  �
  %  W  �  �  �  ,  ]  �  �  �  -  `  �  �  �  *  ]  �  �  �  ,  \  �  �  �  �  �  �    9  _  �  �  �    )  L  u  �  �    =  f  �  �  �  "  \  �  �  �  
	  D	  z	  �	  �	  
  8
  n
  �
  �
    0  `  �  �     0  ^  �  �  �  1  b  �  �  �  ,  V  �  �  �     7  G  K  K  �    7  W  q  �  �  �    2  Q  s  �  �  �  /  Y  �  �  �    M  t  �  �   	  4	  b	  �	  �	  �	  
  8
  f
  �
  �
  �
  "  a  �  �  �  $  S  �  �  �     P    �  �    J  v  �  �  �  �  �  �  �    '  B  [  w  �  �  �    7  T  �  �  �    <  r  �  �  �    J  u  �  �  �  	  C	  x	  �	  �	  �	  
  U
  �
  �
  �
    D  y  �  �    9  k  �  �    =  j  �  �  	  =  B  B  �  �  �  �  �  �    !  <  u  �  �  �  �  #  E  e  �  �  �  �  -  S  l  �  �  �  /  U  u  �  �  	  M	  {	  �	  �	  �	  =
  p
  �
  �
  �
  -  e  �  �  �  '  Q  �  �  �    D  u  �  �  �  �  |    �  �  �  �  �  	  -  S  m  |  �  �  �  �    3  I  f  �  �    /  M  �  �  �    :  `    �  �  	  =	  e	  �	  �	  �	   
  [
  �
  �
  �
    ?  z  �  �  �  0  l  �  �    ,  [  d  F  <  I  j  �  �  �  �  �    +  9  G  [  h  �  �    "  5  U  m  �  �  �  �  !  @  Q  e  �  �  &  H  d  �  �  	  L	  s	  �	  �	  �	  A
  {
  �
  �
  �
  0  q  �  �  �  )  d  �  �    H        :  v  �  �  �  �  �    #  7  J  p  �  �  �  �  �    +  >  W  c  s  �  �  2  T  n  �  �  &  V  v  �  �  	  T	  �	  �	  �	  
  F
  �
  �
  �
  �
  6  y  �  �  	  1  i  �  �  E    �      M  �  �  �  �  �  �  �        C  �  �  �  �  �    a  �  �  �  �    [  �  �  �  �  7  u  �  �  �  (	  e	  �	  �	  �	  "
  Y
  �
  �
  �
  "  N  �  �  �  (  O  ~  �  �  G  *      +  M  z  �  �  �  �  �    2  B  W  _  �  �    &  7  \  �  �  �    0  e  �  �  �    M  �  �  �  	  :	  k	  �	  �	  
  4
  [
  �
  �
    6  \  �  �  �  0  ^  �  �  �    "  V  1  �  8    Y  �  �  �  �  �    j  �  �  �  �    F  p  �  �  �    J  t  �  �  �  0  a  �  �  �  	  T	  �	  �	  �	  
  U
  �
  �
  �
    H    �  �    @  w  �  �    8  v  �  �  6  s  !  L  9  k  �  �    !  '  N  �  �  �    5  f  �  �  �    H  �  �  �  
  6  j  �  �  	  6	  h	  �	  �	  �	  +
  W
  �
  �
  �
  (  V  �  �  �  #  P  �  �  �    N  }  �  �    �    ]  r  �  �  �  �  
  :  a  �  �  �    C  j  �  �    9  e  �  �  �  *  U    �  �  	  J	  u	  �	  �	  
  C
  q
  �
  �
    ?  m  �  �  �  5  i  �  �  �  ,  ^  �  �  �  $  [  �  �  �  J  �  �  �  �  #  C  k  �  �    ;  m  �  �  �  /  b  �  �  �     V  �  �  �  	  L	  ~	  �	  �	  
  A
  x
  �
  �
    ?  t  �  �    :  n  �  �  �  0  d  �  �    6  h  �  �     �    g  �  �    %  i  �  �    +  R  �  �  �    C  w  �  �    <  r  �  �  �  0	  g	  �	  �	  
  2
  f
  �
  �
    0  b  �  �  �  /  `  �  �  �  3  f  �  �     5  i  �  �    7  l  �  C  �  �  �    3  y  �  �    G  w  �  �  !  R  ~  �  �    S  �  �  �  	  Q	  �	  �	  �	  
  N
  �
  �
  �
    M  �  �  �    L  ~  �  �    R  �  �  �     W  �  �  �  $  Z  �  �  Q  r  �  �  �  =  �  �  �    S  �  �    8  l  �  �    Q  �  �  �  4	  k	  �	  �	  
  G
  
  �
  �
  #  X  �  �    :  n  �  �    8  k  �  �    7  h  �  �    6  h  �  �    :  m    �  �  �    c  �  �    E  �  �  �  6  r  �  �  &  _  �  �  	  J	  �	  �	  �	  1
  n
  �
  �
    U  �  �    ;  v  �  �  %  ^  �  �    9  o  �  �    A  v  �  �  �  /  d  �  �  �     �  �    0  �  �  �  #  j  �  �    V  �  �  
  F  }  �  �  8	  s	  �	  �	  #
  b
  �
  �
    O  �  �  �  9  w  �  �  '  a  �  �    M  �  �  �  9  q  �  �  #  _  �  �    H  �  �  �      :  x  �  �    5  v  �  	  3  e  �  �  $  [  �  �  	  C	  {	  �	  �	  #
  a
  �
  �
    D  �  �  �  )  d  �  �    J  �  �  �  2  k  �  �    S  �  �     :  s  �  �     ]  �  7      S  �  �    @  �  �  �  -  Z  |  �  �  @  t  �  �  	  X	  �	  �	  �	  1
  n
  �
  �
    H  �  �  �  )  `  �  �    C  {  �  �  '  ]  �  �    A  x  �  �  "  [  �  �    ?  z    U  �  �    $  (  G  �  �  )  N  u  �  �  6  k  �  �  	  M	  �	  �	  �	  #
  ^
  �
  �
    6  m  �  �    K  �  �  �  +  a  �  �    ?  v  �  �    U  �  �  �  2  j  �  �    J  �    A  �  �    9  o  �  �    H  a  �  �    V  |  �  �  /	  k	  �	  �	  
  C
  �
  �
  �
    X  �  �    5  m  �  �    L  �  �  �  +  b  �  �    ?  v  �  �    S  �  �  �  3  j  �    '  (  )  /  :  u  �  (  M  g  �  �  "  e  �  �  �  !	  f	  �	  �	  �	  )
  j
  �
  �
    7  v  �  �    L  �  �  �  0  b  �  �    E  x  �  �     X  �  �  �  1  k  �  �    E  ~  �  +  1  3  K  P  b  �    ;  X  |  �    Q  {  �  �  (	  h	  �	  �	  �	  6
  u
  �
  �
    F  �  �  �  (  [  �  �  �  1  g  �  �  	  A  x  �  �    M  �  �  �  #  Z  �  �  �  2  h  �  �  .      6    �  �  "  W  u  �  �  0  g  �  �  �  7	  z	  �	  �	  �	  K
  �
  �
  �
    ^  �  �  	  7  q  �  �  "  S  �  �  �  5  i  �  �    G  |  �  �    V  �  �  �  4  j  �  �    3      D  �  �    >  Y  �  �    M  t  �  �  	  W	  �	  �	  �	  
  X
  �
  �
  �
  !  a  �  �  
  6  o  �  �  "  N  �  �  �  7  g  �  �    I  }  �  �    Z  �  �  �  1  k  �  �      �  $  c  �  �    0  j  �  �    J  {  �  �  1	  a	  �	  �	  
  @
  u
  �
  �
    M  �  �  �  $  ]  �  �    9  p  �  �    O  �  �  �  &  ^  �  �  �  3  l  �  �    A  z  �  �    �  �    S  �  �  �  5  m  �  �  #  T  �  �  	  B	  t	  �	  �	  )
  `
  �
  �
    D  ~  �  �    ]  �  �    ;  w  �  �     X  �  �    =  u  �  �  "  Y  �  �    <  t  �  �    W  �  �  �    S  �  �    7  r  �  �  (  ]  �  �  	  K	  }	  �	  �	  9
  m
  �
  �
    S  �  �  �  0  o  �  �    N  �  �  �  2  m  �  �    Q  �  �    ;  r  �  �    Y  �  �    <  w  �  �  �    e  �  �    2  p  �  �  #  O  �  �  	  ;	  j	  �	  �	  
  N
  �
  �
  �
  +  f  �  �    >  z  �  �  $  ]  �  �    =  u  �  �     W  �  �    9  p  �  �    ^  �  �    @  y    =  l  �  �    R  �  �  �  .  h  �  �  	  D	  ~	  �	  �	  
  Z
  �
  �
  �
  5  q  �  �    N  �  �  �  .  g  �  �    K  �  �  �  +  c  �  �    E  |  �  �  %  ]  �  �    <  r  �  �  .  `  �  �  	  @  m  �  �    Q  �  �  �  8	  l	  �	  �	  
  N
  �
  �
  �
  1  j  �  �    K  �  �  �  )  c  �  �    @  z  �  �  !  W  �  �    6  j  �  �    G  �  �  �    :  A  �  $  W  �  �  �  #  N  �  �  �  6  g  �  �  	  G	  z	  �	  �	  
  O
  �
  �
  �
     W  �  �  �  0  f  �  �    @  t  �  �    O  �  �  �  )  ]  �  �  �  4  j  �  �    >  u    �  �  �    6  P  �  �    /  [  �  �    9  j  �  �  	  @	  s	  �	  �	  
  =
  u
  �
  �
  
  ?  y  �  �  
  >  w  �  �  	  ?  ~  �  �    E    �  �    L  �  �  �    R  �  �  �  �  �  �  �  �    -  e  �  �    2  Y  �  �  �  .  ^  �  �  �  #	  M	  t	  �	  �	  
  A
  i
  �
  �
  	  ;  g  �  �  �  *  [  �  �  �  !  ]  �  �  �  '  `  �  �  �  '  ]  �  �  �    5  :  ;  ;  �  �  �    3  Z  �  �  �  $  C  o  �  �  �    N  v  �  �  �  /	  g	  �	  �	  �	  
  H
  z
  �
  �
    .  ]  �  �  	  9  g  �  �  �  /  a  �  �  �  %  Z  �  �  �    R  �  �  �  �  �  s  �  �  �    (  J  y  �  �  �    3  Z  }  �  �  �  '  \  �  �  �  �  )	  a	  �	  �	  �	  
  Q
  �
  �
  �
    >  y  �  �    :  l  �  �  
  ;  i  �  �    +  [  �  �  �    &  )  )  I  i  �  �  �  �  �    A  c  {  �  �  �  �  -  V    �  �    B  f  �  �  �  $	  N	  z	  �	  �	  �	  
  O
  �
  �
  �
    C  }  �  �    7  h  �  �    6  a  �  �  �  /  [  �  �  �  �  	    R  }  �  �  �  �  �      ;  T  i  �  �  
  %  E  v  �  �  �    B  o  �  �  �  �  6	  n	  �	  �	  �	  
  M
  �
  �
  �
    =  t  �  �    3  g  �  �  
  7  e  �  �    8  =  =        O  \  b  o  �  �  �  �    (  >  c  �  �  �  �  �    <  e  }  �  �    >  `    �  �  ,	  `	  �	  �	  �	  
  A
  p
  �
  �
    5  h  �  �  �  %  Q  �  �  �    G  ~  �  �  �  �  �  �  '  <  A  J  a  u  �  �  �  �    #  D  `  r  �  �  �  �  *  N  b  �  �  �  �  ,  T  s  �  �  �   	  Q	  u	  �	  �	   
  A
  w
  �
  �
  �
  (  f  �  �  �    W  �  �  �  "  P  �  �  �  �    -  ,  4  F  [  s  �  �  �  �    '  X  o  �  �  �  �  �    *  L  ]  u  �  �  �  �  <  l  �  �  �  (	  e	  �	  �	  �	  
  V
  �
  �
  �
    K  �  �  �    D  |  �  �  !  I  �  �  �  �      $  /  @  O  �  �  �  �       $  4  B  Q  r  �  �  �  �    5  x  �  �  �    ?  ~  �  �  �  #	  c	  �	  �	  �	  $
  T
  �
  �
  �
  $  M    �  �  *  U  ~  �  �  (  W  �  �  �  �  �    (  .  6  Z  �  �  �  �  �  �    @  X  l    �  �    <  X  r  �  �    :  X  }  �  �  	  F	  s	  �	  �	  
  >
  f
  �
  �
    6  a  �  �  �  .  a  �  �  �    Y  �  �  �  �  �  �      >  &  U  ?  �  �  �  �  
    K  �  �  �  �    N  �  �  �  �  %  \  �  �  �  	  ?	  s	  �	  �	  �	  %
  ]
  �
  �
  �
    E  �  �  �  
  8  m  �  �    1  `  �  �  �  �  �  �      =  {  b  �  }  �  �    >  O  b  �  �    %  C  e  �  �  �  $  N  }  �  �  	  @	  j	  �	  �	  	
  G
  r
  �
  �
    =  j  �  �    7  f  �  �  �  0  `  �  �  �  0  d  �  �    �    �  #  l  �  �  �  �    F  y  �  �  �    O  }  �  �    9  i  �  �  �  #	  X	  �	  �	  �	  "
  V
  �
  �
  �
    E  }  �  �    A  w  �  �    9  n  �  �    4  g  �  �  z  �    
  <  3  J  �  �  �  !  K  r  �  �  �    M  �  �  �    @  u  �  �  	  1	  f	  �	  �	  �	  )
  W
  �
  �
  �
  %  U  �  �  �     P  �  �  �    M  |  �  �    E  u  �  �    G  k  �    /  \  �  �  �  �  $  L  t  �  �     R  z  �  �    A  l  �  �  	  7	  h	  �	  �	  �	  -
  \
  �
  �
  �
  *  \  �  �  �  '  Z  �  �  �  "  P  �  �  �    M  �  �  �    Q  �  �  �  �    9  p  �  �    <  l  �  �  �  2  ]  �  �  �  (  Y  �  �  �  $	  U	  �	  �	  �	  
  M
  �
  �
  �
    M  �  �  �    I  }  �  �    F  z  �  �    L    �  �    O  �  �  �    �  �  $  L  �  �  �  !  Y  �  �  �  '  `  �  �  �  ,  ^  �  �  �  .	  a	  �	  �	  �	  .
  b
  �
  �
  �
  ,  a  �  �  �  ,  `  �  �  �  ,  _  �  �     3  e  �  �    9  l  �  �  
  ?  r  �  
  C  \  �  �    X  �  �  �  ,  i  �  �    @  {  �  �  	  U	  �	  �	  
  8
  n
  �
  �
    L  �  �  �  )  `  �  �    <  u  �  �    K  ~  �  �    E  {  �  �    G  }  �  �    �  _  X  �  �  �  1  o  �  �    W  �  �    @  }  �  �  $	  \	  �	  �	  
  E
  z
  �
  �
  -  d  �  �    I  �  �  �  )  d  �  �    E    �  �  +  b  �  �    I  |  �  �    B  u  �  �  p  �  �  �    Y  �  �    :  v  �  �    K  �  �   	  6	  p	  �	  �	  !
  Z
  �
  �
    ?  z  �  �  #  a  �  �    G  �  �  �  /  g  �  �    P  �  �  �  7  p  �  �    W  �  �    �  �  �  �    E  �  �  �    R  �  �  �  3  p  �  �  	  S	  �	  �	  
  :
  p
  �
  �
    T  �  �  �  2  l  �  �    K  �  �  �  1  h  �  �    L  �  �  �  ,  d  �  �    E  ~  �  �  �  �  �  �  W  �  �  �  #  S  �  �  �    R  �  �  	  6	  n	  �	  �	  
  P
  �
  �
  �
  3  h  �  �    G    �  �  $  _  �  �    =  v  �  �    V  �  �  �  5  l  �  �    K  �  �  �  �  �  8  s  �  �  �  �  5  �  �  �    S  �  �  	  3	  n	  �	  �	  
  M
  �
  �
  �
  *  `  �  �     <  t  �  �    N  �  �  �  +  b  �  �  	  ?  t  �  �    Q  �  �  �  ,  c  �  �    �  �  a  �  �  �    A    �  �    0  o  �  �  	  H	  �	  �	  
  3
  f
  �
  �
    M  �  �  �  *  d  �  �    ?  x  �  �    U  �  �  �  2  i  �  �    C  z  �  �    S  �  �  �  .  �  �  �  �  �  �    y  �  �    B  �  �  �  !	  N	  {	  �	  �	  +
  Y
  �
  �
  �
  :  k  �  �    I    �  �    X  �  �  �  0  j  �  �    D  }  �  �  $  Y  �  �    8  n  �  �    L  �  �  �  �  �    T  �  �  �  -  _  �  �  	  >	  y	  �	  �	  
  I
  �
  �
  �
     V  �  �  �  0  g  �  �    =  t  �  �    O  �  �  �  +  _  �  �    ;  p  �  �    K  �  �  �  $  [  �  {  �  �  �    U  �  �  �  2  s  �  �  	  F	  �	  �	  �	  &
  `
  �
  �
    >  v  �  �    R  �  �  �  0  f  �  �    D  y  �  �    V  �  �  �  1  h  �  �  
  A  z  �  �    V  �  �  f  y  �  �  6  r  �  �  �  2  v  �  �  	  >	  �	  �	  �	  
  Q
  �
  �
    5  i  �  �    M  �  �  �  /  c  �  �    A  x  �  �    T  �  �  �  .  f  �  �    A  y  �  �    U  �  �  M  �  �    1  i  �  �    A  y  �  �  	  O	  �	  �	  �	  $
  ]
  �
  �
    :  o  �  �    P  �  �  �  2  g  �  �    F  }  �  �    U  �  �  �  .  e  �  �  
  @  v  �  �    R  �  ;  K  �  �  �  '  c  �  �    G  �  �  �  &	  d	  �	  �	  
  B
  �
  �
  �
  %  _  �  �    D  {  �  �  *  `  �  �    E  |  �  �  '  a  �  �    A  {  �  �  #  [  �  �    >  v  �  �  ,  R  {  �  �  6  n  �  �    M  �  �  �  .	  n	  �	  �	  
  P
  �
  �
  �
  3  l  �  �    O  �  �     8  n  �  �    U  �  �  �  :  r  �  �    Y  �  �     :  v  �  �    W  �  �      T  w  �  �  1  e  �  �    C  {  �  �  	  Y	  �	  �	  �	  .
  j
  �
  �
    E  �  �  �  *  _  �  �  	  @  |  �  �  &  ]  �  �    <  t  �  �    S  �  �  �  1  l  �  �    U  �  �  �  �  �  %  [  �  �     3  c  �  �  	  D	  u	  �	  �	  
  P
  �
  �
  �
    X  �  �  �  0  h  �  �    9  p  �  �    J  �  �  �  #  X  �  �  �  3  g  �  �    A  u  �  �    H  l  v  p  �  �    5  h  �  �    =  m  �  �  	  G	  {	  �	  �	  
  J
  |
  �
  �
  &  W  �  �  �  -  `  �  �  �  1  k  �  �    ;  s  �  �    I  �  �  �    R  �  �  �  &  c  �  �  �  �  �  Z  �  �  �    E  v  �  �    <  k  �  �  �  0	  l	  �	  �	  
  2
  o
  �
  �
    ;  o  �  �  
  ;  l  �  �    J  {  �  �    K    �  �    H  {  �  �    N  �  �  �      !  !  !  ;  v  �  �  �    B  k  �  �  �  (  X  �  �  �  	  E	  �	  �	  �	  
  2
  k
  �
  �
    -  ^  �  �    3  a  �  �  �  /  a  �  �  �  /  a  �  �  �  3  f  �  �  �  .  `  z  �  �  �  �    9  _  �  �  �  �  .  W  ~  �  �  �  .  _  �  �  �  	  T	  �	  �	  �	   
  7
  i
  �
  �
  �
  #  P  y  �  �    4  g  �  �     :  r  �  �    ?  q  �  �  �  2  h  �  �  �          �    9  W  s  �  �  �    8  V  x  �  �    4  W  �  �  �  	  2	  g	  �	  �	  �	  
  +
  _
  �
  �
  �
    ?  �  �  �    J  x  �  �    C  o  �  �  	  >  n  �  �    5  h  �  �  �  �  �  �    )  B  X  p  �  �  �    +  P  t  �  �  �    ,  Z  �  �  �  �  	  Y	  �	  �	  �	  
  K
  �
  �
  �
    6  p  �  �    .  c  �  �  �  (  Z  �  �  �    J  |  �  �  
    "  "  �  �  �  �    1  G  i  �  �  �  �  �    +  O  s  �  �  �  '  R  o  �  �  �  %	  M	  w	  �	  �	  �	  
  O
  
  �
  �
  �
  <  z  �  �  	  3  d  �  �    2  ^  �  �  �  1  \  �  �  �  �  �  �  �  �      *  :  _  ~  �  �  �  �  �  %  R  l  �  �  �  �    4  W  �  �  �  �  	  J	  }	  �	  �	  �	  0
  i
  �
  �
  �
  #  \  �  �  �    Q  �  �  �  #  P  �  �  �  &  R  W  W  s    �  �  �  �      F  h  y  �  �  �  �      5  K  n  �  �  �  �  �  !  W  �  �  �  �  =	  e	  �	  �	  �	  
  C
  f
  �
  �
  �
     ]  �  �  �    H  {  �  �    ;  o  �  �    0  b  i  ~  �  �  �  �    4  P  ]  m  {  �  �  �  �    (  C  i  �  �  �  �    4  O  j  �  �  �  �  �  +	  j	  �	  �	  �	  
  W
  �
  �
  �
    G  �  �  �    B  w  �  �    F  t  �  �  T  Z  i  �  �  �  �      4  P  b  q  �  �  �      +  A  U  f  �  �  �  �  �    (  C  r  �  �   	  	  H	  �	  �	  �	  
  9
  k
  �
  �
    ;  e  �  �    ?  h  �  �    =  m  �  �  ^  g  y  �  �  �  �  �  �  "  E  Q  ^  x  �  �  �  �  �  
  /  V  q  �  �  �  �  (  Z  {  �  �  �  7	  a	  �	  �	  �	  
  L
  w
  �
  �
    ;  l  �  �  �  *  `  �  �  �  $  [  �  �  �  r  b  s  w  �  �  �  �    !  ;  D  T  ^  x  �  �  �  
  !  3  V  �  �  �    &  Z  �  �  �  	  8	  m	  �	  �	  �	  *
  ^
  �
  �
  �
    K  �  �  �    <  p  �  �    8  g  �  �    5  �  z  s  �  �  �  �  �  �  !    R  �  �  �  �  �    B  n  �  �  �  
  >  ^  }  �  �  	  ;	  d	  �	  �	  �	  (
  Q
  |
  �
  �
    E  n  �  �  �  7  k  �  �  �  &  ]  �  �  �    N  �  �  �  �  �  �  �  �  $    6  /  P  �  �  �  �    C    �  �  �    M  �  �  �  	  5	  j	  �	  �	  �	  "
  U
  �
  �
  �
  (  Z  �  �  �    N  �  �  �    J  }  �  �    E  u  �  �    e  �  �  �  �  �  �     G  g  ~  �  �  �  /  V  x  �  �  �  *  U  �  �  �  	  F	  s	  �	  �	  	
  E
  q
  �
  �
    9  g  �  �  �  0  b  �  �  �  ,  ]  �  �  �  #  W  �  �  �    O  �  F  �  �  �  �  �  �  A  m  �  �  �    K  t  �  �  �  :  f  �  �  �  '	  X	  �	  �	  �	  
  M
  ~
  �
  �
  
  <  s  �  �    ;  p  �  �    5  h  �  �  �  0  b  �  �  �  )  \  �  �  �  -  q  �  �  #  =  B  u  �  �  �  '  e  �  �  �  *  Z  �  �  �  	  L	  �	  �	  �	  
  I
  
  �
  �
  
  ;  p  �  �    <  p  �  �  	  :  l  �  �     2  d  �  �  �  3  h  �  �    4  d  -  v  �  �  )  Z  �  �  �    @  {  �  �     1  d  �  �  �  .	  a	  �	  �	  �	  -
  \
  �
  �
  �
  .  _  �  �  �  ,  ^  �  �  �  *  \  �  �  �  (  Z  �  �  �  .  `  �  �  �  1  d  �  �  G  �  �    0  d  �  �    >  o  �  �    ?  p  �  �  	  <	  p	  �	  �	  
  <
  q
  �
  �
  
  =  q  �  �  
  =  q  �  �  
  =  q  �  �  
  ?  w  �  �    D  z  �  �    K    �  �    �  �  �    E  x  �    9  f  �  �    M  ~  �  �  	  ^	  �	  �	  �	  4
  r
  �
  �
    E  �  �  �  (  [  �  �    =  q  �  �    Q  �  �  �  '  Z  �  �  �  #  X  �  �  �  %  Z  �  �  �     %  A  `  �  �    O  t  �  �  >  r  �  �  	  \	  �	  �	  �	  7
  x
  �
  �
    T  �  �    :  p  �  �  "  V  �  �     ;  q  �  �    R  �  �  �  .  i  �  �    C  x  �  �    H  q  I  P  \  y  �    @  k  �  �  !  [  �  �  �  +	  l	  �	  �	  
  N
  �
  �
  �
  ,  d  �  �    D  z  �  �  +  a  �  �    A  x  �  �    X  �  �  �  6  o  �  �    N  �  �  �  /  h  d  [  v  �  �  �  >  k  �  �  �  O  y  �  �  	  Z	  �	  �	  �	  0
  q
  �
  �
    J  �  �  �  -  b  �  �    C  x  �  �    V  �  �  �  2  j  �  �    F  ~  �  �  #  Y  �  �    <  t  �  ^  b  �    F  f  �  �     9  z  �  �  �  7	  �	  �	  �	  
  K
  �
  �
  �
  (  `  �  �    A  u  �  �  &  Y  �  �    <  q  �  �    N  �  �  �  (  a  �  �    <  s  �  �    Q  �  l  �  �  -  b  |  �  �  �  9  x  �  �  �  @	  ~	  �	  �	  
  R
  �
  �
  �
  '  ]  �  �  
  ;  m  �  �    Q  �  �  �  &  _  �  �  �  6  o  �  �    E    �  �  !  V  �  �  �  3  h  �  \  �    M  l  }  �  �    T  �  �  �  	  _	  �	  �	  �	  &
  q
  �
  �
    @  �  �  �  '  Y  �  �  
  =  q  �  �    N  �  �  �  )  _  �  �    8  o  �  �    H  ~  �  �  #  [  �  �    �  z  D  V  �  �    K  u  �  �  		  L	  �	  �	  �	  
  G
  �
  �
  �
    T  �  �  
  5  g  �  �     N  ~  �  �  3  f  �  �    D  z  �  �    T  �  �  �  ,  e  �  �  
  @  x  �  �  �  /  8  *  e  �  �    K  v  �  �  )	  ]	  �	  �	  �	  /
  j
  �
  �
    ;  v  �  �    L  �  �  �  -  `  �  �    @  t  �  �    S  �  �  �  (  b  �  �    8  q  �  �    J  �  �  �  �      3  d  �  �    L  �  �   	  :	  l	  �	  �	  
  P
  �
  �
  �
  "  _  �  �     5  o  �  �    I    �  �  ,  `  �  �    @  v  �  �    R  �  �  �  +  c  �  �  
  B  x  �  �     m  �    C  x  �     3  W  �  �  	  ?	  m	  �	  �	  
  O
  �
  �
  �
    _  �  �  �  1  n  �  �    F    �  �  (  [  �  �    =  q  �  �    Q  �  �  �  *  c  �  �    =  u  �  �      �    M  �  �  �  2  b  �  �  	  F	  x	  �	  �	  
  V
  �
  �
  �
  )  e  �  �    :  u  �  �    M  �  �  �  .  b  �  �    C  x  �  �    T  �  �  �  +  d  �  �    ;  t  �  �    �  �     M  �  �  �  9  g  �  �  	  M	  �	  �	  �	  (
  d
  �
  �
    A  |  �  �     Y  �  �    ;  t  �  �    V  �  �    :  q  �  �    U  �  �  �  5  o  �  �    N  �  �  �  /  g  �  �    M  �  �  �  /  b  �  �  	  I	  	  �	  �	  /
  f
  �
  �
    L  �  �  �  (  f  �  �    D  ~  �  �  *  a  �  �    F  }  �  �  %  _  �  �  	  B  |  �  �  $  \  �  �    >  w  �  �    8  l  �  �    Q  �  �  �  2	  j	  �	  �	  
  F
  {
  �
  �
    U  �  �    6  o  �  �    H    �  �  .  c  �  �  
  @  u  �  �    R  �  �  �  ,  c  �  �    L  �  �  �    �    >  p  �  �    N  |  �  �  	  V	  �	  �	  �	  &
  _
  �
  �
  �
  *  _  �  �    5  h  �  �    6  i  �  �    =  r  �  �    B  v  �  �    I  }  �  �    O  �  �  �          �  �  -  Y  �  �  �  &  Y  �  �  �  	  Q	  �	  �	  �	  
  R
  }
  �
  �
    L  z  �  �    C  r  �  �  �  /  j  �  �  �  0  f  �  �    7  l  �  �    6  i  �  �    A  d  u  y  y  z  �  �    C  `  �  �  �  $  J  r  �  �  	  &	  U	  �	  �	  �	  
  B
  �
  �
  �
    7  b  �  �  �    G  }  �  �  ,  [  �  �  �     T  �  �  �    K    �  �    S  �  �  �  �  �  �  �  �  �  �    3  U  �  �  �  �    L  s  �  �  �  	  I	  �	  �	  �	  �	  
  T
  �
  �
  �
    D  }  �  �    C  t  �  �    D  o  �  �    =  n  �  �    C  o  �  �    5  W  h  k  k  l  u  �  �  �      B  m  �  �  �  �    9  f  �  �  �  	  P	  {	  �	  �	  �	  -
  \
  �
  �
  �
    9  c  �  �  �    M  �  �  �  %  ]  �  �  �  (  Y  �  �  �    P  �  �  �  �  �  �  �  Y  �  �  �  �  �  
  -  Q  j  �  �  �  �  /  R  n  �  �  �  		  4	  f	  �	  �	  �	  �	  !
  V
  �
  �
  �
  
  9  {  �  �    A  s  �  �    =  j  �  �    ;  j  �  �    5  f  �  �  �  �  I  w  �  �  �  �  �    (  P  g  |  �  �  �  �    6  V  z  �  �  �  	  =	  q	  �	  �	  �	  ,
  e
  �
  �
  �
    O  }  �  �    :  o  �  �  �  -  _  �  �  �  %  S  �  �  �    8  <  <  <  e  �  �  �  �  �  �  	  ,  ?  R  l  �  �  �  �  �    A  s  �  �  �  	  )	  I	  s	  �	  �	  �	  
  /
  i
  �
  �
  �
    Y  �  �  �  %  S  �  �  �  $  P    �  �  !  S    �  �  �  �  .  P  v  |  �  �  �  �  �    %  =  Q  u  �  �  �  �    )  H  c    �  �  �  �  	  -	  b	  �	  �	  �	  
  F
  ~
  �
  �
  
  ;  r  �  �    8  i  �  �    <  h  �  �    >  l  �  �  �  +  D  g  r  z  �  �  �  �      6  O  j  �  �  �  �  �       9  V  p  �  �  �  	  *	  V	  �	  �	  �	  �	  
  (
  U
  �
  �
  �
  	  :  u  �  �    4  g  �  �    5  c  �  �    6  e  �  $  2  N  g  u  �  �  �  �  �      5  C  e  �  �  �  �  �    E  ^  x  �  �  �  �  	  #	  :	  S	  p	  �	  �	  
  *
  K
  w
  �
  �
    >  g  �  �    ?  k  �  �    :  k  �  �  �  4  k    "  :  a  t  �  �  �  �  �      ,  =  _  �  �  �  �  �      .  C  e  �  �  �  �  �  &	  b	  �	  �	  �	  
  :
  m
  �
  �
  �
    W  �  �  �    G  �  �  �    =  r  �  �  
  9  l    )  6  ]  k  �  �  �  �  �         >  [  i  x  �  �  �  �    #  :  V  w  �  �  	  +	  O	  ~	  �	  �	  
  4
  ^
  �
  �
     )  W  �  �  �    G  w  �  �    ?  t  �  �    A  o  �     )  D  S  p  �  �  �  �  �  �      (  @  P  �  �  �  �  �    E  |  �  �  �  	  N	  |	  �	  �	  �	  $
  W
  �
  �
  �
    K  y  �  �    ;  l  �  �  �  )  b  �  �  �    T  �  �  �  2  3  9  O  Q  �  �  �  �  �  �    <  8  \  e  �  �  �  "  0  S  �  �  �  	  2	  _	  �	  �	  �	  
  F
  y
  �
  �
    1  a  �  �  �  !  P  �  �  �    G  w  �  �    B  m  �  �    7  2  S  9  X  l  x  �  �  �  �  �    G  u  �  �  �  �  5  d  �  �  �  �  0	  [	  �	  �	  �	  
  K
  x
  �
  �
    :  n  �  �    A  r  �  �    6  k  �  �  �  1  f  �  �  �  *  ^  �  �    Q  \  8  s  J  �  �       ,  :  p  �  �    '  K  w  �  �  	  1	  e	  �	  �	  �	  $
  T
  �
  �
  �
  !  R  �  �  �    F  v  �  �    A  t  �  �    <  n  �  �    :  j  �  �    1  �  8  l  T  �  �  �  �  $  S    �  �  �    I  z  �  �  	  =	  o	  �	  �	  
  2
  `
  �
  �
  �
  +  X  �  �  �    R  �  �  �    P  ~  �  �    I  |  �  �    E  t  �  �    ?  s  �  �  &  f  �  �  �  �    N  x  �  �    C  p  �  �  	  4	  e	  �	  �	  �	  *
  \
  �
  �
  �
  )  U  �  �  �    N  �  �  �    N  �  �  �    L    �  �    C  w  �  �    I  {  �  �    �  #  h  �  �  	  0  o  �  �  �    N  �  �  �  	  F	  {	  �	  �	  	
  B
  w
  �
  �
    8  n  �  �  	  :  o  �  �    8  l  �  �    7  j  �  �    ;  q  �  �  
  >  t  �  �    B  w  �  .  p  �  �    2  q  �  �    H  x  �  �  	  H	  |	  �	  �	  
  I
  ~
  �
  �
    J  ~  �  �    K  }  �  �    M  ~  �  �    M    �  �     T  �  �  �  #  Y  �  �  �  '  ]  �  �  1  U  �  �  �    W  �  �    8  m  �  �  	  M	  �	  �	  �	  2
  d
  �
  �
    G  }  �  �    U  �  �  �  ,  e  �  �    @  w  �  �     U  �  �  �  (  R  �  �  �  #  T  �  �  �  !  S  E  �  �  �    >  w  �  �    L  �  �  	  =	  q	  �	  �	  *
  ^
  �
  �
    D  z  �  �  $  ^  �  �    :  r  �  �    Q  �  �  �  5  k  �  �    N  �  �  �    R  �  �  �    G  z  �  %  �  �    '  e  �  �    H    �  �  %	  S	  �	  �	  
  >
  p
  �
  �
    Z  �  �  �  2  m  �  �    E  �  �  �  )  `  �  �  
  @  w  �  �    V  �  �  �  3  k  �  �    B  t  �  �      *  5  m  �  �    -  X  �  �  	  E	  v	  �	  �	  /
  `
  �
  �
    E  z  �  �  !  Z  �  �  �  1  j  �  �    F  }  �  �  $  [  �  �    8  o  �  �    I  �  �  �  #  V  �  �  �  S      D  �  �  
  4  g  �  �  	  ;	  d	  �	  �	  
  N
  z
  �
  �
  ,  c  �  �  �  :  v  �  �    K  �  �  �  &  ^  �  �  
  =  u  �  �    T  �  �  �  1  f  �  �    9  k  �  �  �    J  �  �      &  F  �  �  	  6	  d	  �	  �	  
  E
  v
  �
  �
    N  �  �  �    Y  �  �  �  .  h  �  �    A  w  �  �    S  �  �  �  3  h  �  �    E  {  �  �    V  �  �  �      4  �  �  �  �     Z  �  �  �  3	  q	  �	  �	  
  I
  �
  �
  �
  -  `  �  �    ?  s  �  �    P  �  �  �  +  a  �  �    <  r  �  �    N  �  �  �  (  _  �  �    8  p  �  �      (  5  $  �  �  �  )  v  �  �  	  6	  {	  �	  �	   
  O
  �
  �
  	  :  j  �  �    Q  �  �  �  .  e  �  �    ?  x  �  �    R  �  �  �  -  d  �  �    A  x  �  �    T  �  �  �        �  �  �  �    I  |  �  �  	  K	  �	  �	  �	  (
  [
  �
  �
    ?  o  �  �    T  �  �  �  1  i  �  �    B  |  �  �    U  �  �  �  1  g  �  �    D  z  �  �     V  �  �  �        t  �  �  �    G  �  �  �  $	  a	  �	  �	  
  =
  u
  �
  �
  #  U  �  �     9  m  �  �    M  �  �  �  $  a  �  �    :  u  �  �    O  �  �  �  /  e  �  �    D  {  �  �  
  
  
  �  [  �  �  �    Y  �  �  �  '	  b	  �	  �	  
  :
  s
  �
  �
    P  �  �  �  3  g  �  �    G  }  �  �     Z  �  �  �  3  m  �  �    G  �  �  �  '  \  �  �    <  r  �  �  �  �  �  z  A  y  �  �  "  Z  �  �  �  /	  i	  �	  �	  
  >
  x
  �
  �
    O  �  �  �  .  b  �  �  
  A  w  �  �    T  �  �  �  0  h  �  �  
  A  y  �  �    S  �  �  �  0  e  �  �        (  ?  v  �  �    R  �  �  �  .	  i	  �	  �	  
  E
  �
  �
  �
  $  ^  �  �    :  u  �  �    T  �  �  �  5  k  �  �    N  �  �  �  -  d  �  �    F  }  �  �  %  ]  �  �            A  u  �  �    J    �  �  (	  a	  �	  �	  
  F
  ~
  �
  �
    \  �  �    :  r  �  �    T  �  �  �  3  k  �  �    H  �  �  �  )  ^  �  �    <  q  �  �    Q  �  �  �  �  �  �  �  ,  \  �  �    :  i  �  �  	  J	  ~	  �	  �	   
  [
  �
  �
  �
  0  h  �  �    G  ~  �  �  "  U  �  �  �  :  n  �  �    G  |  �  �    S  �  �  �  '  ]  �  �    ?  t  �  �  �  �  A  m  �  �  �    N  �  �  �  	  7	  l	  �	  �	  �	  /
  b
  �
  �
    $  R  �  �  �  +  U  �  �  �  /  [  �  �  �  0  b  �  �  �  )  _  �  �  �  (  b  �  �  �  *  ]  �  �  �  �  �  �  3  ]  �  �  �  �    M  {  �  �  �  &	  Z	  �	  �	  �	  
  Q
  �
  �
  �
    ;  s  �  �    0  Z  �  �  �    I  y  �  �    H  �  �  �    M  �  �  �    C  w  �  �    3  D  G  G  I  $  K  i  �  �  �  �  !  M  m  �  �  �   	  E	  i	  �	  �	  �	  
  F
  �
  �
  �
    %  I  y  �  �    0  d  �  �    E  s  �  �    <  m  �  �  �  2  g  �  �  �  8  l  �  �  �  �  �  �    6  J  g  �  �  �  �    ;  O  y  �  �  �  	  2	  W	  �	  �	  �	  �	  
  Q
  �
  �
  �
    A  |  �  �    <  q  �  �  
  8  f  �  �  �  .  ^  �  �     2  `  �  �  �  (  P  b  f  e  g  �    6  U  m  �  �  �  �      2  R  v  �  �  �  	  ;	  n	  �	  �	  �	  
  <
  c
  �
  �
  �
    4  b  �  �  �    K  �  �  �  '  ^  �  �  �  ,  [  �  �  �    T  �  �  �  �  �  �  �  �    /  H  ^  q  �  �  �  �  �  	  +  Y  �  �  �  �  	  "	  @	  d	  �	  �	  �	  �	  
  =
  s
  �
  �
  �
  '  Z  �  �  �  ,  ^  �  �  �  *  X  �  �  �  )  X  �  �  �  &  X  �  �  �  �  �  �    )  <  P  a  �  �  �  �  �    '  C  ^  u  �  �  �  �  	  	  4	  c	  �	  �	  �	  
  ?
  w
  �
  �
  �
    J  ~  �  �  �  +  a  �  �  �  (  V  �  �  �  $  R  �  �  �  "  O  r  z  z  �  �     2  C  W  z  �  �  �  �  �  �  &  E  \  r  �  �  �  	  	  3	  [	  ~	  �	  �	  �	  �	  
  2
  U
  �
  �
  �
    ;  m  �  �    B  r  �  �    A  n  �  �    <  m  �  �    5  ?  ?  �  �    ,  6  P  d  �  �  �  �  �  �    E  ^  u  �  �  �  �  �  	  7	  Q	  k	  �	  �	  �	  �	  $
  G
  m
  �
  �
    3  \  �  �  �    O  �  �  �    D  w  �  �    @  q  �  �        �  �    *  /  K  T  v  �  �  �  �  �    0  D  Y  i  �  �  �  �  �  	  ?	  r	  �	  �	  �	  �	  
  6
  W
  y
  �
  �
  �
    G  k  �  �    5  ^  �  �  �  *  ]  �  �  �  "  W  �  �  �    �  �  �     -  D  N  m  �  �  �  �  �  �    7  P  c  }  �  �  �  
	   	  :	  Q	  q	  �	  �	  �	  �	  �	  
  O
  �
  �
  �
  �
  .  b  �  �  �    N  �  �  �    @  u  �  �    9  l  �  �    �  �  �    /  @  L  i  ~  �  �  �  �  �    =  N  m  �  �  �  �  �  �  	  5	  M	  f	  �	  �	  �	  
  ?
  `
  �
  �
  �
  !  L  p  �  �    <  h  �  �  �  6  c  �  �  �  &  Y  �  �  �     �  �  �    -  B  I  h  p  �  �  �  �  �    '  5  J  b  p  �  �  �  �  	  ,	  a	  �	  �	  �	  
  8
  p
  �
  �
  �
    H  �  �  �    A  u  �  �  �  /  c  �  �  �  )  \  �  �  �  #  R  �  �  �       B  R  d  z  �  �  �  �  �  �    7  X  j  �  �  �  �  2	  R	  k	  �	  �	   
  ,
  Q
  w
  �
  �
  	  5  a  �  �  �  +  V  �  �  �    L  y  �  �    G  t  �  �  
  ?  n  �  �  �  �       A  W  X  r  �  �  �  �  �      5  r  �  �  �  	  :	  n	  �	  �	  �	  
  D
  s
  �
  �
  �
  ,  ]  �  �  �    J  z  �  �    4  i  �  �  �  *  \  �  �  �     Q  �  �  �  �    �      ,  \    d  �  �  �  �  *  N  Y  x  �  �  	  1	  W	  �	  �	  �	  

  6
  g
  �
  �
  �
  &  U  �  �  �    Z  �  �  �  !  R  �  �  �    L  }  �  �    H  x  �  �    J  |  �  	  	  �  &  �  A  �  �  �  �  �  !  ]  �  �  �  �  !	  U	  �	  �	  �	  
  B
  o
  �
  �
  �
  0  a  �  �  �  2  b  �  �  �  #  V  �  �  �  !  U  �  �  �    O  �  �  �    J  }  �  �  �  �  $  �  4  6  ]  �  �  �  -  L  h  �  �  �  %	  W	  �	  �	  �	  
  E
  y
  �
  �
  	  9  n  �  �    1  b  �  �  �  ,  _  �  �  �  (  Z  �  �  �  &  W  �  �  �    P  �  �  �    S  �  �    M  ~  �  �  �  �    S  �  �  �  	  E	  t	  �	  �	  
  <
  h
  �
  �
    6  f  �  �  �  -  \  �  �  �  +  ]  �  �  �  *  \  �  �  �  '  T  �  �  �     S  �  �  �    Q  �  �  ~  �    G  w  �  �    ;  [  �  �  �  +	  T	  �	  �	  �	  "
  R
  ~
  �
  �
    P  ~  �  �    J    �  �    K  }  �  �    H  |  �  �    F  z  �  �    L  �  �  �    H  y  �  �    �  �    S    �  �    \  �  �  �  	  ]	  �	  �	  �	  
  U
  �
  �
  �
  "  V  �  �  �  %  X  �  �  �  %  X  �  �  �  &  Y  �  �  �  '  Y  �  �  �  .  `  �  �  �  (  [  �  �  �  "  T  �  �  D  x  �  �  �  F  �  �  �  	  R	  �	  �	  �	  (
  a
  �
  �
    ?  v  �  �  '  V  �  �  �    G  u  �  �    9  h  �  �  �  /  _  �  �  �  %  V  �  �  �    P  �  �  �    I  {    K  x  �  �  �    k  �  �  �  /	  �	  �	  �	  
  P
  �
  �
    5  m  �  �    G  q  �  �    ,  X  �  �  �    G  u  �  �  	  ;  k  �  �  �  /  _  �  �  �  "  U  �  �  �    P  �  �  �  �  �  �    Z  �  �  �  #	  f	  �	  �	  �	  .
  k
  �
  �
    G  �  �  �    8  i  �  �  �    B  q  �  �  �  /  `  �  �  �  &  V  �  �  �    L    �  �    G  w  �  �    B  t  �  �  �  �    =  �  �  �  �  A	  �	  �	  �	  
  V
  �
  �
  
  6  n  �  �    5  M  i  �  �  �    8  h  �  �  �  &  U  �  �  �    I  y  �  �    B  t  �  �    ;  l  �  �    3  e  �  �  �  �  f  �  �  �  �  -	  n	  �	  �	  �	  .
  o
  �
  �
    D  �  �     0  R  t  �  �  �    0  W  �  �  �    1  _  �  �  �     R  �  �  �    H  |  �  �    C  u  �  �    =  m  �  �  -  |  �    �  �  	  Q	  �	  �	  �	  
  X
  �
  �
  �
  (  _  �  �    =  p  �  �  �    5  ]  �  �  �    5  c  �  �  �    M  |  �  �    @  r  �  �    7  i  �  �  �  0  b  �  �  �  g  f  h  p  �  �  #	  V	  �	  �	  �	  /
  l
  �
  �
    >  {  �  �    O  x  �  �  �  -  \  �  �  �    ?  l  �  �  �  &  T  �  �  �    E  w  �  �    =  o  �  �    4  e  m  m  �  �  �  ;  [  �  �  �  7	  l	  �	  �	   
  B
  }
  �
  �
    Q  �  �  �  (  a  �  �  �    5  b  �  �  �    E  w  �  �    8  j  �  �  �  0  c  �  �  �  ,  ^  �  �  �  &  W  l  l  l  x  -  5  (  `  �  �  	  @	  s	  �	  �	  
  L
  �
  �
  �
    Z  �  �  �  0  i  �  �    '  P  ~  �  �    1  `  �  �  �    L  |  �  �    B  t  �  �  	  ;  m  �  �    5  d  |  |  |  r  �    8  h  �  �  	  E	  	  �	  �	  
  [
  �
  �
  �
  3  p  �  �    I  �  �  �    I  s  �  �  �  $  R  �  �  �  
  :  i  �  �     2  d  �  �  �  +  ]  �  �  �  #  R  f  o  o  o  6  �     7  g  �  �  	  I	  ~	  �	  �	  
  Y
  �
  �
  �
  0  j  �  �    D  }  �  �  !  M  y  �  �    /  ^  �  �  �    M  ~  �  �    D  v  �  �    ?  p  �  �  	  :  \  b  b  b  b  �  �  �  &  ^  �  �  �  6	  m	  �	  �	  
  G
  }
  �
  �
    V  �  �  �  0  g  �  �    A  v  �  �  �  ,  Z  �  �  �    I  |  �  �    C  u  �  �    >  p  �  �    7  \  i  i  i  i  �  �  �    R  �  �  �  ,	  _	  �	  �	  �	  9
  l
  �
  �
    E  {  �  �    U  �  �  �  ,  d  �  �     1  `  �  �  �    J  {  �  �    A  v  �  �    >  q  �  �    6  T  c  d  d  d  n  �  �    <  l  �  �  	  ?	  q	  �	  �	  
  M
  �
  �
  �
  "  S  �  �  �  2  d  �  �    <  r  �  �    E  {  �  �    H  y  �  �    A  s  �  �    >  q  �  �    4  K  R  S  S  S  Q  �  �  �    L  ~  �  �  	  C	  x	  �	  �	  
  A
  z
  �
  �
    K  �  �  �  (  `  �  �  �  *  [  �  �  �  <  q  �  �    ;  q  �  �    =  p  �  �    >  t  �  �    H  R  R  R  R  �  �    .  I  j  �  �  �  	  /	  \	  �	  �	  �	  
  ;
  g
  �
  �
  �
    @  x  �  �    ?  p  �  �    E  n  �  �    K  x  �  �    @  p  �  �    B  t  �  �    7  o  �  �  �  �  �  �  �  �    (  I  o  �  �  �  �  	  E	  s	  �	  �	  �	  
  W
  �
  �
  �
  �
  7  l  �  �  �    H  s  �  �  �  6  d  �  �    :  n  �  �    <  o  �  �  �  .  c  �  �  �  !  3  6  7  9  �  �  �  �    ,  V  z  �  �  �  �  	  P	  u	  �	  �	  �	  
  .
  T
  �
  �
  �
    "  F  w  �  �    .  d  �  �    A  p  �  �  
  <  l  �  �    6  h  �  �  �  :  n  �  �  �  �  �  �  �  �  �  �       C  f  �  �  �  �  �  	  4	  S	  t	  �	  �	  �	  �	  
  B
  z
  �
  �
  �
  ,  e  �  �  �  #  T  �  �  �    B  v  �  �    ;  i  �  �    @  o  �  �    ;  d  |  �  �  �  �  �  �  �  �    4  W  t  �  �  �  �  �  	  '	  F	  j	  �	  �	  �	  �	  (
  R
  t
  �
  �
  �
    1  W  �  �  �    >  p  �  �    J  �  �  �    O  }  �  �    F  z  �  �    *  0  2  2  �  �  �  �  �    )  N  h  z  �  �  �  �  	  *	  E	  b	  �	  �	  �	  �	  �	  
  3
  N
  n
  �
  �
  �
    H  y  �  �    C  v  �  �    B  q  �  �    @  q  �  �    <  p  �  �  �  �  �  �  �  �  �  �  �  �  $  N  d  y  �  �  �  �  �  	  !	  F	  f	  �	  �	  �	  �	  
  0
  Q
  p
  �
  �
  �
    *  N  t  �  �    ,  V  �  �  �  %  Q    �  �    O  ~  �  �    L  }  �  �  �  �  �  �  �  �  �  �     A  V  g  �  �  �  �  �  �  	  9	  `	  �	  �	  �	  �	  �	  
  5
  T
  r
  �
  �
  �
  �
  "  O  x  �  �  �  0  e  �  �  �  (  [  �  �  �    T  �  �  �    N  �  �  �  �  �  �  �  �  �  �    .  O  b  x  �  �  �  �  �  	  9	  R	  m	  �	  �	  �	  �	  �	  
  *
  K
  w
  �
  �
  �
    N    �  �     *  U  ~  �  �    =  n  �  �    7  h  �  �  �  0  ]  �  �  �  �  �  �  �  �  �     %  P  c  q  �  �  �  �  �  	  	  :	  [	  v	  �	  �	  �	  �	  '
  K
  k
  �
  �
  �
  �
  �
    @  n  �  �  �    K  }  �  �    1  i  �  �    3  b  �  �  �  +  Z  �  �  �  �  �  �  �  �  �    G  Z  h  �  �  �  �  �  �  	  ,	  U	  �	  �	  �	  �	  �	  �	  
  @
  ^
  t
  �
  �
  �
    =  b  �  �  �    H  t  �  �    :  j  �  �  �  +  `  �  �  �     X  �  �  �  �  �  �  �  �  �    6  O  m  {  �  �  �  �  �   	  9	  O	  g	  x	  �	  �	  �	  �	  �	  
  4
  a
  �
  �
  �
    A  t  �  �     &  U  �  �  �    M    �  �    E  v  �  �    >  p  �  �  �  �  �  �  �  �  �    #  G  j  �  �  �  �  �  �  �  	  )	  O	  o	  �	  �	  �	  �	  
  M
  q
  �
  �
  �
  "  P  w  �  �  �  7  d  �  �  �  )  W  �  �  �    I  x  �  �    G  x  �  �    �  �  �  �  �  �      ,  G  h  v  �  �  �  �  �  
	  	  3	  E	  v	  �	  �	   
  
  F
  |
  �
  �
    )  Y  �  �  �    I  ~  �  �    6  l  �  �  �  +  \  �  �  �  &  U  �  �  �     P  �  �  �  �  �  �    	  (  5  K  w  �  �  �  �  �  &	  X	  }	  �	  �	  �	  
  K
  n
  �
  �
  �
  "  K  y  �  �    8  c  �  �  �  )  U  �  �  �    L  {  �  �    ?  r  �  �    5  f  �  �  �  �  �  �  �  	  /    D  8  g  �  �  �  	  '	  ^	  �	  �	  �	  
  .
  Z
  �
  �
  �
    D  u  �  �     0  b  �  �    5  i  �  �  �  .  _  �  �  �  (  Z  �  �  �  #  U  �  �  �  '  �  �  �  �  �  �  �  4  Y  m  �  �  �  	  /	  Z	  	  �	  �	   
  -
  Z
  �
  �
  �
    E  t  �  �  
  E  s  �  �    <  k  �  �  �  3  d  �  �  �  0  `  �  �  �  (  [  �  �  �  #  U  �  o  �  �  �  �  �    E  t  �  �  �  	  C	  o	  �	  �	  �	  5
  a
  �
  �
  �
    T  �  �  �    H  y  �  �    6  l  �  �    5  i  �  �  �  ,  ^  �  �  �  &  X  �  �  �    S  �  �  �  E  �  �  �  "  ,  /  k  �  �  �  $	  \	  �	  �	  �	  
  L
  �
  �
  �
  	  <  q  �  �    4  g  �  �  �  %  X  �  �  �    M  ~  �  �    D  u  �  �    <  l  �  �    4  f  �  �  �  -  .  r  �  �    S  }  �  �  	  *	  b	  �	  �	  
  *
  Y
  �
  �
  �
    F  p  �  �    2  ^  �  �  �  $  R  �  �  �    D  t  �  �    9  i  �  �  �  .  _  �  �  �  #  V  �  �  �    M  =  v  �  �  %  W  }  �  �  1	  c	  �	  �	  �	  
  5
  \
  �
  �
  �
    B  o  �  �    .  Z  �  �  �    L  z  �  �    @  n  �  �     1  a  �  �  �  %  V  �  �  �    R  �  �  �    J  y  �  �     F  i  �  �  %	  T	  �	  �	  �	  �	  
  
  G
  {
  �
  �
    .  Z  �  �  �    ?  n  �  �  �  *  Y  �  �  �  "  Q  �  �  �    G  v  �  �    ?  o  �  �    6  j  �  �     4  �  �    T  c  �  �  	  F	  l	  �	  �	  �	  
  -
  M
  d
  �
  �
  �
  �
    B  p  �  �  �    E  t  �  �  �  1  g  �  �  �  &  W  �  �  �    O  �  �  �    D  u  �  �    D  v  �  �    �  l  `  S  x  �  	  9	  b	  �	  �	  
  !
  7
  N
  e
  �
  �
  �
  �
  �
    ,  G  f  �  �  �  &  S  �  �  �    <  m  �  �    5  f  �  �  �  ,  ^  �  �  �  &  X  �  �  �    N  �  �  �  �  a  s  �  �  �  <	  O	  p	  �	  �	  �	  
  5
  h
  �
  �
  �
  �
  �
    0  O  u  �  �  �  �  "  T  �  �  �     .  a  �  �  �    P  �  �  �    K  }  �  �    C  t  �  �    ;  m  �  �  �  c  e  �  	   	  &	  3	  k	  �	  �	  
  9
  Q
  m
  �
  �
  �
    '  C  a  |  �  �  �  �  &  I  f  �  �  �    >  k  �  �  �  ,  Z  �  �  �    Q  �  �  �    I  {  �  �    C  u  �  �  s  �  �  	  I	  �  	  ?	  }	  �	  �	  +
  N
  k
  �
  �
  �
  �
  �
    9  [  �  �  �    *  L  p  �  �  �    C  p  �  �  �  $  R  �  �  �    C  v  �  �  
  :  m  �  �    5  g  �  �  �  a  {  	  �  �  �  	  K	  �	  �	  �	  /
  _
  �
  �
  �
  �
  �
    1  T  v  �  �  �    <  m  �  �  �    I  w  �  �  �  +  Z  �  �  �    G  y  �  �    @  r  �  �    :  l  �  �  �  �  �  	  	  �  �  �  %	  ^	  �	  �	  	
  :
  n
  �
  �
  �
  �
    2  P  q  �  �  �  �  !  D  i  �  �  �    N  {  �  �    =  l  �  �    4  f  �  �  �  .  `  �  �  �  (  Z  �  �  �  �  �  �  �  �  �  �  �  .	  f	  �	  �	  
  <
  t
  �
  �
  �
  �
    :  \  �  �  �  �    <  _  �  �  �    :  g  �  �  �    M  ~  �  �    A  s  �  �  	  :  l  �  �    5  g  �  �  �  �  �  �  M  b  �  �  �  -	  e	  �	  �	  
  D
  {
  �
  �
  �
  �
    7  ]  �  �  �     (  S  �  �  �     +  Y  �  �  �    ;  j  �  �  �  .  _  �  �  �  (  X  �  �  �  "  T  �  �  �  �  �  �  �  .  S  �  �  �  +	  e	  �	  �	  
  @
  x
  �
  �
  �
       @  e  �  �  �  �  )  V  �  �  �    2  `  �  �  �    L  |  �  �    ?  q  �  �    9  l  �  �    6  i  �  �  �  �  �  �  B    G  y  �  �  	  Y	  �	  �	  �	  )
  d
  �
  �
  �
    -  O  s  �  �  �    ,  Q  x  �  �     .  \  �  �  �    F  v  �  �  
  ;  m  �  �    6  i  �  �     2  e  �  �  �  �  �  �  �  	  ?  n  �  �  	  >	  v	  �	  �	  
  E
  }
  �
  �
    -  N  t  �  �  �    4  ^  �  �  �    1  _  �  �  �    D  t  �  �  	  9  k  �  �    9  k  �  �    6  g  �  �  �  �  �  �  �    5  c  �  �  �   	  V	  �	  �	  �	  
  O
  �
  �
  �
    =  d  �  �  �    .  ]  �  �  �    1  ^  �  �  �    F  v  �  �    =  o  �  �  	  <  p  �  �    ;  m  �  �  �  �  �  �  �  �  !  J  j  �  �  �  &	  Q	  u	  �	  �	  
  1
  c
  �
  �
  �
  ,  X  �  �  �  #  N  x  �  �  �    K  x  �  �  	  :  k  �  �    7  j  �  �    5  h  �  �    4  g  �  �  �  �  �  �  C  f  �  �  �  �  �  %	  G	  c	  |	  �	  �	  �	  
  2
  ]
  �
  �
  �
  �
    H  u  �  �  �    O  |  �  �    I  z  �  �    K  �  �  �    P  �  �  �  !  V  �  �  �  (  Y  z  �  �  �  �  F  i  |  �  �  �  �  	  .	  A	  Y	  y	  �	  �	  �	  
  &
  N
  �
  �
  �
  �
    S  �  �  �     &  M  w  �  �    <  i  �  �    D  u  �  �    C  v  �  �    7  l  �  �  	  .  B  F  G  I  H  d  m  }  �  �  �  	   	  3	  M	  n	  �	  �	  �	  �	  
  8
  X
  v
  �
  �
  �
    +  I  n  �  �  �  (  T  �  �  �  .  _  �  �  �  .  ^  �  �  �  (  \  �  �  �  $  _  �  �  �  �  �  �  �  H  _  g  x  �  �  �  	  	  .	  G	  k	  �	  �	  �	  �	  �	  
  0
  J
  e
  
  �
  �
    ,  R  �  �  �    2  [  �  �  �    B  p  �  �    @  l  �  �  	  B  s  �  �    =  q  �  �  �  �  �  L  a  i  |  �  �  �  �  	  	  3	  V	  |	  �	  �	  �	  �	  
  7
  W
  o
  �
  �
  �
  �
    2  Q  o  �  �  �    E  n  �  �    <  k  �  �    9  k  �  �  �  1  e  �  �  �  .  `  �  �  �  �  Q  m  q  �  �  �  �  �  		  	  1	  W	  	  �	  �	  �	  �	   
  
  7
  Q
  q
  �
  �
  �
  �
    3  ^  �  �  �    8  h  �  �  �  %  T  �  �  �    I  z  �  �    C  u  �  �  	  9  _  k  m  m  K  l  y  �  �  �  �  �  	  	  <	  ]	  v	  �	  �	  �	  �	  �	  
  $
  ?
  _
  �
  �
  �
  �
    ?  ^  |  �  �  �    <  j  �  �  �    L    �  �  	  >  s  �  �    7  k  �  �    .  \  h  h  E  i  y  �  �  �  �  �  �  	  ,	  ?	  a	  �	  �	  �	  �	  �	  
  7
  P
  h
  �
  �
  �
  �
       1  M  p  �  �  �  $  L  z  �  �    5  c  �  �  �  .  ^  �  �  �  '  W  �  �  �  "  V  `  `  7  d  }  �  �  �  �  �  �  	  '	  7	  \	  �	  �	  �	  �	  �	   
  
  3
  J
  k
  �
  �
  �
  �
  �
  ,  Z  �  �  �    )  S  ~  �  �     ,  [  �  �  �    F  z  �  �    B  t  �  �    7  i  k  7  e    �  �  �  �  �  �  	   	  ?	  d	  }	  �	  �	  �	  �	  �	  
  %
  ;
  Y
  
  �
  �
  �
    9  U  n  �  �  �  �  %  W  }  �  �    4  c  �  �  �     T  �  �  �    J  }  �  �    ?  v  9  Z  u  �  �  �  �  �  �  	  	  5	  Q	  a	  �	  �	  �	  �	  �	  

  6
  V
  n
  �
  �
  �
  �
  �
    $  =  ]  �  �  �    ?  l  �  �  �  (  P  �  �  �    K  {  �  �    C  q  �  �    @  q  A  Q  i  �  �  �  �  �  �  	   	  .	  G	  Y	  ~	  �	  �	  �	  �	  
  
  0
  G
  _
  
  �
  �
  �
  �
    O  �  �  �  �  (  Y  �  �  �  
  @  t  �  �    4  g  �  �  �  +  ]  �  �  �  $  X  �  :  L  R  �  �  �  �  �  �  	   	  7	  E	  f	  �	  �	  �	  �	  �	  �	  
  #
  6
  M
  i
  �
  �
  �
    ?  m  �  �     '  N  }  �  �    @  s  �  �    4  b  �  �  �  )  W  �  �  �  )  Y  �  �  8  I  V  s  �  �  �  �  �  �  	  +	  9	  O	  c	  }	  �	  �	  �	  �	  �	  (
  a
  �
  �
  �
  �
  +  ^  �  �  �  	  8  g  �  �  �  +  [  �  �  �    N  }  �  �    A  w  �  �    8  l  �  �     w  �    R  h  �  �  �  �  �  	  %	  J	  D	  h	  n	  �	  �	   
  %
  >
  d
  �
  �
  �
    D  q  �  �  �  '  W  �  �  �    ?  o  �  �    .  _  �  �  �  )  U  �  �  �    P  |  �  �    F  �  �  �  1  q  �  �  �  �  �  �  	  T	  �	  �	  �	  �	  
  <
  f
  �
  �
  �
    4  _  �  �  �    J  w  �  �    8  l  �  �    ?  p  �  �    4  h  �  �  �  0  c  �  �  �  )  \  �  �  �  �  �  0  \  [  �  �  �  	  $	  <	  s	  �	  �	  �	  
  ?
  k
  �
  �
  �
  '  X  �  �  �    B  t  �  �    <  p  �  �  �  .  _  �  �  �  '  Y  �  �  �     P  �  �  �    J  |  �  �    �      =  K  w  �  �  	  9	  _	  v	  �	  �	   
  '
  Q
  ~
  �
  �
    ;  g  �  �  �  '  S  �  �  �    >  m  �  �    3  b  �  �  �  *  Y  �  �  �    R  �  �  �    J  |  �  �    E  �  '  8  '  3  X  t  �  �  *	  B	  i	  �	  �	  �	   
  D
  l
  �
  �
    .  [  �  �  �    L  |  �  �    ?  m  �  �    2  a  �  �  �  &  V  �  �  �    O  �  �  �    G  z  �  �    @  �      C  t  �  �  �  �  �  	  %	  _	  �	  �	  �	  
  C
  p
  �
  �
    3  _  �  �  �  $  R  �  �  �    F  u  �  �  
  :  i  �  �  �  0  `  �  �  �  ,  ]  �  �  �  $  X  �  �  �    �    N  \  u  �  �  �  �  �  �  	  B	  k	  �	  �	  �	  
  M
  {
  �
  �
  �
  '  X  �  �  �    C  u  �  �    ;  n  �  �    0  a  �  �  �  %  U  �  �  �  #  S  �  �  �  "  S  �  �  �    H  t  �  �  �  �  �  �  �  	  ,	  F	  `	  �	  �	  �	  �	  /
  R
  q
  �
  �
  �
  )  T  �  �  �    E  q  �  �    6  j  �  �  �  /  b  �  �  �  #  U  �  �  �    O  �  �  �    M  �  �  O  _  �  �  �  �  �  �  �  	  3	  G	  `	  y	  �	  �	  �	  �	  �	  
  9
  l
  �
  �
  �
  %  R  �  �  �    ;  l  �  �    3  c  �  �  �  ,  ]  �  �  �  "  R  �  �  �    K  �  �  �    N  �  a  p    �  �  �  �  �  �  &	  N	  k	  �	  �	  �	  �	  �	  �	  
  D
  [
  v
  �
  �
  �
    D  n  �  �  �    L  z  �  �  	  ;  p  �  �    3  d  �  �  �  *  ^  �  �  �  %  V  �  �  �  "  U  w  x  �  �  �  �  �  	  	  3	  M	  m	  �	  �	  �	  �	  
  %
  ?
  \
  z
  �
  �
  �
  �
    1  P  y  �  �    :  g  �  �  �  *  W  �  �  �    N    �  �    J  |  �  �    C  u  �  �  	  <  |  y  �  �  �  �  �  	  -	  F	  a	  �	  �	  �	  �	  �	  
  &
  W
  �
  �
  �
  �
  �
    ;  _  �  �  �  �    P    �  �  �  -  b  �  �  �  !  T  �  �  �    M  �  �  �    G  y  �  �    @  v  �  �  �  �  �  	  1	  I	  b	  x	  �	  �	  �	  �	  
  
  ;
  _
  �
  �
  �
  �
  -  Q  m  �  �  �  �  #  M  y  �  �  �  0  \  �  �  �    H  v  �  �    ?  q  �  �    7  i  �  �  �  1  V  w  �  �  �  �  �  	  5	  S	  t	  �	  �	  �	  �	  �	  
  8
  V
  u
  �
  �
  �
  �
    >  d  �  �  �  (  R    �  �    4  a  �  �  �    I  y  �  �    @  q  �  �    9  l  �  �  �  0  :  :  u  �  �  �  �  �  	  9	  X	  {	  �	  �	  �	  �	  
  *
  R
  s
  �
  �
  �
  �
    1  W    �  �  �  %  U  �  �  �    <  o  �  �  �  0  c  �  �  �  +  ]  �  �  �  '  X  �  �  �     4  4  4  z  �  �  �  �  	   	  ?	  ]	  }	  �	  �	  �	  �	  
  ,
  Y
  
  �
  �
  �
    1  T  y  �  �  �    ?  m  �  �  �  "  O  {  �  �    ?  o  �  �    6  h  �  �  �  0  c  �  �  �  (  B  B  B  y  �  �  �  �  	  ,	  I	  b	  ~	  �	  �	  �	  �	  

  1
  [
  �
  �
  �
  �
    ;  ^  �  �  �    4  ]  �  �  �    ?  k  �  �  �  '  Y  �  �  �     S  �  �  �    N  �  �  �    &  0  0  0  y  �  �  �  �  	  <	  V	  p	  �	  �	  �	  �	   
  !
  D
  f
  �
  �
  �
  �
    4  Y  �  �  �    7  c  �  �  �    H  w  �  �    7  i  �  �  �  1  c  �  �  �  .  `  �  �  �    !  !  !  !  t  }  �  �  �  	  6	  T	  t	  �	  �	  �	  �	  
  +
  O
  p
  �
  �
  �
  �
    @  e  �  �  �    0  _  �  �  �    @  n  �  �    5  f  �  �  �  1  d  �  �  �  /  b  �  �  �    (  (  (  (  d  x  �  �  �  	  ,	  J	  k	  �	  �	  �	  �	  �	  
  B
  n
  �
  �
  �
    *  L  p  �  �  �    7  d  �  �  �    L  x  �  �    =  q  �  �    A  u  �  �  
  >  s  �  �  �    &  &  &  &  R  s  �  �  �  �  "	  D	  c	  	  �	  �	  �	  �	  
  5
  a
  �
  �
  �
  �
  '  H  f  �  �  �    7  c  �  �  �  $  W  �  �  �    N  �  �  �    Q  �  �  �  !  T  �  �  �    '  ,  -  -  -  D  i  �  �  �  �  	  :	  e	  �	  �	  �	  �	  �	  
  @
  g
  �
  �
  �
  �
    A  b  �  �  �    2  ^  �  �  �  *  Y  �  �  �  ,  ^  �  �  �  /  `  �  �  �  /  f  �  �  �  -  J  Q  Q  Q  Q  